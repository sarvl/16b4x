LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

USE work.p_arithmetic.to_uint;
USE work.p_mem.t_mem_rbyte;

ENTITY flash_data IS
	PORT(
		clk      : IN    std_ulogic;

		addr     : IN    std_ulogic_vector(22 DOWNTO 0);
		data_in  : IN    std_ulogic_vector(15 DOWNTO 0);
		data_out :   OUT std_ulogic_vector(15 DOWNTO 0);
		we       : IN    std_ulogic
	);
END ENTITY;


ARCHITECTURE arch OF flash_data IS 
	SIGNAL flash : t_mem_rbyte(65535 * 2 + 1 DOWNTO 0) := (
		00000=>x"A0",00001=>x"0E",00002=>x"48",00003=>x"00",00004=>x"0E",
		00005=>x"06",00006=>x"98",00007=>x"02",00008=>x"29",00009=>x"9A",
		00010=>x"59",00011=>x"2E",00012=>x"A7",00013=>x"1F",00014=>x"58",
		00015=>x"24",00016=>x"A0",00017=>x"20",00018=>x"48",00019=>x"08",
		00020=>x"40",00021=>x"4A",00022=>x"00",00023=>x"4D",00024=>x"C8",
		00025=>x"02",00026=>x"AF",00027=>x"00",00028=>x"2F",00029=>x"A7",
		00030=>x"18",00031=>x"1C",00052=>x"AF",00053=>x"00",00054=>x"AF",
		00055=>x"00",00056=>x"AF",00057=>x"00",00058=>x"AF",00059=>x"00",
		00060=>x"A0",00061=>x"0E",00062=>x"48",00063=>x"00",00064=>x"A1",
		00065=>x"1E",00066=>x"5F",00067=>x"21",00068=>x"A1",00069=>x"3E",
		00070=>x"00",00071=>x"2D",00072=>x"C8",00073=>x"22",00074=>x"C8",
		00075=>x"02",00076=>x"2F",00077=>x"C7",00078=>x"A0",00079=>x"00",
		00080=>x"0F",00081=>x"00",00082=>x"0F",00083=>x"02",00084=>x"A1",
		00085=>x"10",00086=>x"0F",00087=>x"1F",00088=>x"18",00089=>x"26",
		00120=>x"AF",00121=>x"00",00122=>x"AF",00123=>x"00",00124=>x"AF",
		00125=>x"00",00126=>x"AF",00127=>x"00",00128=>x"58",00129=>x"21",
		00130=>x"A0",00131=>x"00",00132=>x"6A",00133=>x"00",00134=>x"A0",
		00135=>x"00",00136=>x"6A",00137=>x"02",00138=>x"6A",00139=>x"04",
		00140=>x"6A",00141=>x"06",00142=>x"A0",00143=>x"02",00144=>x"0F",
		00145=>x"00",00146=>x"A2",00147=>x"00",00148=>x"0F",00149=>x"02",
		00150=>x"A0",00151=>x"02",00152=>x"58",00153=>x"22",00154=>x"68",
		00155=>x"00",00156=>x"A1",00157=>x"F2",00158=>x"48",00159=>x"E0",
		00160=>x"58",00161=>x"2E",00162=>x"5D",00163=>x"19",00174=>x"AF",
		00175=>x"00",00176=>x"A3",00177=>x"12",00178=>x"48",00179=>x"00",
		00180=>x"58",00181=>x"2E",00182=>x"5D",00183=>x"19",00184=>x"A2",
		00185=>x"14",00186=>x"48",00187=>x"00",00188=>x"1F",00189=>x"FB",
		00220=>x"AF",00221=>x"00",00222=>x"AF",00223=>x"00",00224=>x"A0",
		00225=>x"02",00226=>x"48",00227=>x"00",00228=>x"19",00229=>x"2A",
		00440=>x"AF",00441=>x"00",00442=>x"A0",00443=>x"0A",00444=>x"48",
		00445=>x"00",00446=>x"1F",00447=>x"FB",00528=>x"A0",00529=>x"04",
		00530=>x"48",00531=>x"00",00532=>x"19",00533=>x"DA",01004=>x"AF",
		01005=>x"00",01006=>x"AF",01007=>x"00",01008=>x"A0",01009=>x"06",
		01010=>x"48",01011=>x"00",01012=>x"19",01013=>x"FA",01024=>x"58",
		01025=>x"28",01026=>x"58",01027=>x"00",01028=>x"58",01029=>x"28",
		01030=>x"58",01031=>x"10",01512=>x"AF",01513=>x"00",01514=>x"AF",
		01515=>x"00",01516=>x"AF",01517=>x"00",01518=>x"AF",01519=>x"00",
		01520=>x"A0",01521=>x"08",01522=>x"48",01523=>x"00",01524=>x"19",
		01525=>x"FA",01536=>x"58",01537=>x"28",01538=>x"59",01539=>x"08",
		02030=>x"AF",02031=>x"00",02032=>x"A0",02033=>x"0A",02034=>x"48",
		02035=>x"00",02036=>x"19",02037=>x"5A",02048=>x"6F",02049=>x"01",
		02050=>x"58",02051=>x"22",02052=>x"60",02053=>x"06",02054=>x"C0",
		02055=>x"02",02056=>x"58",02057=>x"22",02058=>x"68",02059=>x"06",
		02060=>x"67",02061=>x"01",02062=>x"09",02063=>x"00",02064=>x"6F",
		02065=>x"01",02066=>x"6F",02067=>x"23",02068=>x"0E",02069=>x"18",
		02070=>x"F8",02071=>x"16",02072=>x"00",02073=>x"34",02074=>x"5F",
		02075=>x"21",02076=>x"E0",02077=>x"00",02078=>x"C2",02079=>x"20",
		02080=>x"01",02081=>x"0D",02082=>x"67",02083=>x"01",02084=>x"67",
		02085=>x"23",02086=>x"09",02087=>x"00",02088=>x"A0",02089=>x"20",
		02090=>x"0F",02091=>x"20",02092=>x"0F",02093=>x"20",02094=>x"A1",
		02095=>x"22",02096=>x"0F",02097=>x"3F",02098=>x"58",02099=>x"22",
		02100=>x"60",02101=>x"20",02102=>x"01",02103=>x"54",02104=>x"58",
		02105=>x"22",02106=>x"C0",02107=>x"40",02108=>x"02",02109=>x"0D",
		02110=>x"C0",02111=>x"22",02112=>x"58",02113=>x"22",02114=>x"68",
		02115=>x"20",02116=>x"58",02117=>x"2E",02118=>x"5D",02119=>x"19",
		02380=>x"AF",02381=>x"00",02382=>x"AF",02383=>x"00",02384=>x"A0",
		02385=>x"0C",02386=>x"48",02387=>x"00",02388=>x"18",02389=>x"AA",
		02560=>x"A0",02561=>x"0E",02562=>x"48",02563=>x"00",02564=>x"19",
		02565=>x"FA",03066=>x"AF",03067=>x"00",03068=>x"AF",03069=>x"00",
		03070=>x"AF",03071=>x"00",03072=>x"A0",03073=>x"10",03074=>x"48",
		03075=>x"00",03076=>x"19",03077=>x"AA",03498=>x"AF",03499=>x"00",
		03500=>x"AF",03501=>x"00",03502=>x"AF",03503=>x"00",03504=>x"A0",
		03505=>x"12",03506=>x"48",03507=>x"00",03508=>x"18",03509=>x"3A",
		03520=>x"58",03521=>x"28",03522=>x"A0",03523=>x"00",03524=>x"C8",
		03525=>x"02",03526=>x"2F",03527=>x"E7",03528=>x"AF",03529=>x"00",
		03530=>x"AC",03531=>x"00",03532=>x"02",03533=>x"AA",03534=>x"17",
		03535=>x"F1",03536=>x"48",03537=>x"24",03538=>x"17",03539=>x"ED",
		03540=>x"48",03541=>x"02",03542=>x"17",03543=>x"E9",03544=>x"A0",
		03545=>x"42",03546=>x"48",03547=>x"46",03548=>x"17",03549=>x"E3",
		03550=>x"A0",03551=>x"40",03552=>x"48",03553=>x"46",03554=>x"17",
		03555=>x"DD",03556=>x"05",03557=>x"4B",03558=>x"AC",03559=>x"00",
		03560=>x"AF",03561=>x"00",03562=>x"AF",03563=>x"00",03564=>x"AF",
		03565=>x"00",03566=>x"AF",03567=>x"00",03568=>x"A0",03569=>x"14",
		03570=>x"48",03571=>x"00",03572=>x"19",03573=>x"C2",03574=>x"AF",
		03575=>x"00",03576=>x"AF",03577=>x"00",03578=>x"A1",03579=>x"E6",
		03580=>x"48",03581=>x"E0",03582=>x"1F",03583=>x"FB",03584=>x"A0",
		03585=>x"C0",03586=>x"48",03587=>x"04",03588=>x"48",03589=>x"06",
		03590=>x"A3",03591=>x"10",03592=>x"A0",03593=>x"20",03594=>x"17",
		03595=>x"C1",03596=>x"A6",03597=>x"48",03598=>x"17",03599=>x"B1",
		03600=>x"C8",03601=>x"42",03602=>x"2F",03603=>x"D3",03604=>x"A0",
		03605=>x"62",03606=>x"A3",03607=>x"10",03608=>x"17",03609=>x"B3",
		03610=>x"A0",03611=>x"54",03612=>x"17",03613=>x"A3",03614=>x"C8",
		03615=>x"42",03616=>x"2F",03617=>x"D3",03618=>x"C8",03619=>x"62",
		03620=>x"2F",03621=>x"87",03622=>x"A0",03623=>x"18",03624=>x"17",
		03625=>x"A3",03626=>x"A0",03627=>x"02",03628=>x"17",03629=>x"9F",
		03630=>x"A0",03631=>x"0C",03632=>x"17",03633=>x"9B",03634=>x"A0",
		03635=>x"22",03636=>x"AF",03637=>x"00",03638=>x"A4",03639=>x"10",
		03640=>x"17",03641=>x"93",03642=>x"A4",03643=>x"02",03644=>x"17",
		03645=>x"8F",03646=>x"A4",03647=>x"12",03648=>x"17",03649=>x"8B",
		03650=>x"A4",03651=>x"18",03652=>x"17",03653=>x"87",03654=>x"A2",
		03655=>x"00",03656=>x"17",03657=>x"83",03658=>x"A4",03659=>x"1E",
		03660=>x"17",03661=>x"7F",03662=>x"A4",03663=>x"1A",03664=>x"17",
		03665=>x"7B",03666=>x"A4",03667=>x"1C",03668=>x"17",03669=>x"77",
		03670=>x"A4",03671=>x"12",03672=>x"17",03673=>x"73",03674=>x"A5",
		03675=>x"06",03676=>x"17",03677=>x"6F",03678=>x"A5",03679=>x"06",
		03680=>x"17",03681=>x"6B",03682=>x"A4",03683=>x"12",03684=>x"17",
		03685=>x"67",03686=>x"A4",03687=>x"02",03688=>x"17",03689=>x"63",
		03690=>x"A4",03691=>x"10",03692=>x"17",03693=>x"5F",03694=>x"A1",
		03695=>x"E4",03696=>x"48",03697=>x"E0",03698=>x"0B",03699=>x"00",
		03700=>x"1F",03701=>x"FF",04022=>x"AF",04023=>x"00",04024=>x"A0",
		04025=>x"16",04026=>x"48",04027=>x"00",04028=>x"1F",04029=>x"FB",
		04030=>x"58",04031=>x"22",04032=>x"60",04033=>x"00",04034=>x"0F",
		04035=>x"00",04036=>x"A1",04037=>x"20",04038=>x"A0",04039=>x"42",
		04040=>x"88",04041=>x"04",04042=>x"28",04043=>x"94",04044=>x"88",
		04045=>x"06",04046=>x"28",04047=>x"F4",04048=>x"5F",04049=>x"21",
		04050=>x"A0",04051=>x"02",04052=>x"6A",04053=>x"02",04054=>x"0F",
		04055=>x"3F",04056=>x"0F",04057=>x"5F",04058=>x"58",04059=>x"30",
		04060=>x"58",04061=>x"00",04062=>x"5F",04063=>x"21",04064=>x"A0",
		04065=>x"04",04066=>x"6A",04067=>x"02",04068=>x"0F",04069=>x"3F",
		04070=>x"0F",04071=>x"5F",04072=>x"58",04073=>x"30",04074=>x"58",
		04075=>x"00",04076=>x"AF",04077=>x"00",04078=>x"58",04079=>x"22",
		04080=>x"60",04081=>x"02",04082=>x"58",04083=>x"22",04084=>x"60",
		04085=>x"24",04086=>x"1E",04087=>x"03",04088=>x"AF",04089=>x"00",
		04090=>x"AF",04091=>x"00",04092=>x"AF",04093=>x"00",04094=>x"A0",
		04095=>x"08",04096=>x"0F",04097=>x"1F",04098=>x"A0",04099=>x"00",
		04100=>x"A0",04101=>x"22",04102=>x"A0",04103=>x"EE",04104=>x"88",
		04105=>x"E0",04106=>x"28",04107=>x"6C",04108=>x"AF",04109=>x"00",
		04110=>x"00",04111=>x"54",04112=>x"01",04113=>x"14",04114=>x"02",
		04115=>x"38",04116=>x"C8",04117=>x"E2",04118=>x"2F",04119=>x"B7",
		04120=>x"AF",04121=>x"00",04122=>x"A0",04123=>x"F4",04124=>x"48",
		04125=>x"E0",04126=>x"08",04127=>x"01",08188=>x"AF",08189=>x"00",
		08190=>x"A0",08191=>x"08",08192=>x"0F",08193=>x"1F",08194=>x"A0",
		08195=>x"2E",08196=>x"A0",08197=>x"02",08198=>x"01",08199=>x"10",
		08200=>x"C8",08201=>x"22",08202=>x"2F",08203=>x"D3",08204=>x"A0",
		08205=>x"F8",08206=>x"48",08207=>x"E0",08208=>x"08",08209=>x"01",
		12280=>x"AF",12281=>x"00",12282=>x"AF",12283=>x"00",12284=>x"AF",
		12285=>x"00",
		OTHERS => x"00");
BEGIN
	data_out <= flash(to_uint(addr & '1')) & flash(to_uint(addr & '0'));
	
	PROCESS(ALL) IS BEGIN
		IF rising_edge(clk) THEN
		IF we THEN
			flash(to_uint(addr & '1')) <= data_in(15 DOWNTO 8);
			flash(to_uint(addr & '0')) <= data_in( 7 DOWNTO 0);
		END IF;
		END IF;
	END PROCESS;

END ARCHITECTURE;



LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

USE work.p_arithmetic.to_uint;
USE work.p_mem.t_mem_rword;

ENTITY ram_data IS
	PORT(
		clk   : IN    std_ulogic;

		addr  : IN    std_ulogic_vector(15 DOWNTO 0);
		data  : INOUT std_ulogic_vector(15 DOWNTO 0);
		re    : IN    std_ulogic;
		we    : IN    std_ulogic
	);
END ENTITY;

ARCHITECTURE arch OF ram_data IS 
	--SHOULD contain the same data as flash
	--double check pls
	SIGNAL ram : t_mem_rword(65535 DOWNTO 0) := (
0000=>x"A20E",0001=>x"4800",0002=>x"0E06",0003=>x"9802",0004=>x"299A",
0005=>x"592E",0006=>x"A000",0007=>x"5824",0008=>x"A020",0009=>x"4808",
0010=>x"404A",0011=>x"004D",0012=>x"C802",0013=>x"0111",0014=>x"2FA7",
0015=>x"181C",0016=>x"AF00",0017=>x"AF00",0018=>x"AF00",0019=>x"AF00",
0020=>x"AF00",0021=>x"AF00",0022=>x"AF00",0023=>x"AF00",0024=>x"AF00",
0025=>x"AF00",0026=>x"AF00",0027=>x"AF00",0028=>x"AF00",0029=>x"AF00",
0030=>x"A10E",0031=>x"4800",0032=>x"A11E",0033=>x"5F21",0034=>x"A13E",
0035=>x"002D",0036=>x"C822",0037=>x"C802",0038=>x"2FC7",0039=>x"A000",
0040=>x"0F00",0041=>x"0F02",0042=>x"A110",0043=>x"0F1F",0044=>x"1826",
0045=>x"AF00",0046=>x"AF00",0047=>x"AF00",0048=>x"AF00",0049=>x"AF00",
0050=>x"AF00",0051=>x"AF00",0052=>x"AF00",0053=>x"AF00",0054=>x"AF00",
0055=>x"AF00",0056=>x"AF00",0057=>x"AF00",0058=>x"AF00",0059=>x"AF00",
0060=>x"AF00",0061=>x"AF00",0062=>x"AF00",0063=>x"AF00",0064=>x"5821",
0065=>x"A000",0066=>x"6A00",0067=>x"A000",0068=>x"6A02",0069=>x"6A04",
0070=>x"6A06",0071=>x"A002",0072=>x"0F00",0073=>x"A200",0074=>x"0F02",
0075=>x"A002",0076=>x"5822",0077=>x"6800",0078=>x"A1F2",0079=>x"48E0",
0080=>x"582E",0081=>x"5D13",0082=>x"AF00",0083=>x"AF00",0084=>x"AF00",
0085=>x"AF00",0086=>x"AF00",0087=>x"AF00",0088=>x"A312",0089=>x"4800",
0090=>x"582E",0091=>x"5D13",0092=>x"A214",0093=>x"4800",0094=>x"1FFB",
0095=>x"AF00",0096=>x"AF00",0097=>x"AF00",0098=>x"AF00",0099=>x"AF00",
0100=>x"AF00",0101=>x"AF00",0102=>x"AF00",0103=>x"AF00",0104=>x"AF00",
0105=>x"AF00",0106=>x"AF00",0107=>x"AF00",0108=>x"AF00",0109=>x"AF00",
0110=>x"AF00",0111=>x"AF00",0112=>x"A002",0113=>x"4800",0114=>x"192A",
0115=>x"AF00",0116=>x"AF00",0117=>x"AF00",0118=>x"AF00",0119=>x"AF00",
0120=>x"AF00",0121=>x"AF00",0122=>x"AF00",0123=>x"AF00",0124=>x"AF00",
0125=>x"AF00",0126=>x"AF00",0127=>x"AF00",0128=>x"AF00",0129=>x"AF00",
0130=>x"AF00",0131=>x"AF00",0132=>x"AF00",0133=>x"AF00",0134=>x"AF00",
0135=>x"AF00",0136=>x"AF00",0137=>x"AF00",0138=>x"AF00",0139=>x"AF00",
0140=>x"AF00",0141=>x"AF00",0142=>x"AF00",0143=>x"AF00",0144=>x"AF00",
0145=>x"AF00",0146=>x"AF00",0147=>x"AF00",0148=>x"AF00",0149=>x"AF00",
0150=>x"AF00",0151=>x"AF00",0152=>x"AF00",0153=>x"AF00",0154=>x"AF00",
0155=>x"AF00",0156=>x"AF00",0157=>x"AF00",0158=>x"AF00",0159=>x"AF00",
0160=>x"AF00",0161=>x"AF00",0162=>x"AF00",0163=>x"AF00",0164=>x"AF00",
0165=>x"AF00",0166=>x"AF00",0167=>x"AF00",0168=>x"AF00",0169=>x"AF00",
0170=>x"AF00",0171=>x"AF00",0172=>x"AF00",0173=>x"AF00",0174=>x"AF00",
0175=>x"AF00",0176=>x"AF00",0177=>x"AF00",0178=>x"AF00",0179=>x"AF00",
0180=>x"AF00",0181=>x"AF00",0182=>x"AF00",0183=>x"AF00",0184=>x"AF00",
0185=>x"AF00",0186=>x"AF00",0187=>x"AF00",0188=>x"AF00",0189=>x"AF00",
0190=>x"AF00",0191=>x"AF00",0192=>x"AF00",0193=>x"AF00",0194=>x"AF00",
0195=>x"AF00",0196=>x"AF00",0197=>x"AF00",0198=>x"AF00",0199=>x"AF00",
0200=>x"AF00",0201=>x"AF00",0202=>x"AF00",0203=>x"AF00",0204=>x"AF00",
0205=>x"AF00",0206=>x"AF00",0207=>x"AF00",0208=>x"AF00",0209=>x"AF00",
0210=>x"AF00",0211=>x"AF00",0212=>x"AF00",0213=>x"AF00",0214=>x"AF00",
0215=>x"AF00",0216=>x"AF00",0217=>x"AF00",0218=>x"AF00",0219=>x"AF00",
0220=>x"AF00",0221=>x"A00A",0222=>x"4800",0223=>x"1FFB",0224=>x"AF00",
0225=>x"AF00",0226=>x"AF00",0227=>x"AF00",0228=>x"AF00",0229=>x"AF00",
0230=>x"AF00",0231=>x"AF00",0232=>x"AF00",0233=>x"AF00",0234=>x"AF00",
0235=>x"AF00",0236=>x"AF00",0237=>x"AF00",0238=>x"AF00",0239=>x"AF00",
0240=>x"AF00",0241=>x"AF00",0242=>x"AF00",0243=>x"AF00",0244=>x"AF00",
0245=>x"AF00",0246=>x"AF00",0247=>x"AF00",0248=>x"AF00",0249=>x"AF00",
0250=>x"AF00",0251=>x"AF00",0252=>x"AF00",0253=>x"AF00",0254=>x"AF00",
0255=>x"AF00",0256=>x"AF00",0257=>x"AF00",0258=>x"AF00",0259=>x"AF00",
0260=>x"AF00",0261=>x"AF00",0262=>x"AF00",0263=>x"AF00",0264=>x"A004",
0265=>x"4800",0266=>x"19DA",0267=>x"AF00",0268=>x"AF00",0269=>x"AF00",
0270=>x"AF00",0271=>x"AF00",0272=>x"AF00",0273=>x"AF00",0274=>x"AF00",
0275=>x"AF00",0276=>x"AF00",0277=>x"AF00",0278=>x"AF00",0279=>x"AF00",
0280=>x"AF00",0281=>x"AF00",0282=>x"AF00",0283=>x"AF00",0284=>x"AF00",
0285=>x"AF00",0286=>x"AF00",0287=>x"AF00",0288=>x"AF00",0289=>x"AF00",
0290=>x"AF00",0291=>x"AF00",0292=>x"AF00",0293=>x"AF00",0294=>x"AF00",
0295=>x"AF00",0296=>x"AF00",0297=>x"AF00",0298=>x"AF00",0299=>x"AF00",
0300=>x"AF00",0301=>x"AF00",0302=>x"AF00",0303=>x"AF00",0304=>x"AF00",
0305=>x"AF00",0306=>x"AF00",0307=>x"AF00",0308=>x"AF00",0309=>x"AF00",
0310=>x"AF00",0311=>x"AF00",0312=>x"AF00",0313=>x"AF00",0314=>x"AF00",
0315=>x"AF00",0316=>x"AF00",0317=>x"AF00",0318=>x"AF00",0319=>x"AF00",
0320=>x"AF00",0321=>x"AF00",0322=>x"AF00",0323=>x"AF00",0324=>x"AF00",
0325=>x"AF00",0326=>x"AF00",0327=>x"AF00",0328=>x"AF00",0329=>x"AF00",
0330=>x"AF00",0331=>x"AF00",0332=>x"AF00",0333=>x"AF00",0334=>x"AF00",
0335=>x"AF00",0336=>x"AF00",0337=>x"AF00",0338=>x"AF00",0339=>x"AF00",
0340=>x"AF00",0341=>x"AF00",0342=>x"AF00",0343=>x"AF00",0344=>x"AF00",
0345=>x"AF00",0346=>x"AF00",0347=>x"AF00",0348=>x"AF00",0349=>x"AF00",
0350=>x"AF00",0351=>x"AF00",0352=>x"AF00",0353=>x"AF00",0354=>x"AF00",
0355=>x"AF00",0356=>x"AF00",0357=>x"AF00",0358=>x"AF00",0359=>x"AF00",
0360=>x"AF00",0361=>x"AF00",0362=>x"AF00",0363=>x"AF00",0364=>x"AF00",
0365=>x"AF00",0366=>x"AF00",0367=>x"AF00",0368=>x"AF00",0369=>x"AF00",
0370=>x"AF00",0371=>x"AF00",0372=>x"AF00",0373=>x"AF00",0374=>x"AF00",
0375=>x"AF00",0376=>x"AF00",0377=>x"AF00",0378=>x"AF00",0379=>x"AF00",
0380=>x"AF00",0381=>x"AF00",0382=>x"AF00",0383=>x"AF00",0384=>x"AF00",
0385=>x"AF00",0386=>x"AF00",0387=>x"AF00",0388=>x"AF00",0389=>x"AF00",
0390=>x"AF00",0391=>x"AF00",0392=>x"AF00",0393=>x"AF00",0394=>x"AF00",
0395=>x"AF00",0396=>x"AF00",0397=>x"AF00",0398=>x"AF00",0399=>x"AF00",
0400=>x"AF00",0401=>x"AF00",0402=>x"AF00",0403=>x"AF00",0404=>x"AF00",
0405=>x"AF00",0406=>x"AF00",0407=>x"AF00",0408=>x"AF00",0409=>x"AF00",
0410=>x"AF00",0411=>x"AF00",0412=>x"AF00",0413=>x"AF00",0414=>x"AF00",
0415=>x"AF00",0416=>x"AF00",0417=>x"AF00",0418=>x"AF00",0419=>x"AF00",
0420=>x"AF00",0421=>x"AF00",0422=>x"AF00",0423=>x"AF00",0424=>x"AF00",
0425=>x"AF00",0426=>x"AF00",0427=>x"AF00",0428=>x"AF00",0429=>x"AF00",
0430=>x"AF00",0431=>x"AF00",0432=>x"AF00",0433=>x"AF00",0434=>x"AF00",
0435=>x"AF00",0436=>x"AF00",0437=>x"AF00",0438=>x"AF00",0439=>x"AF00",
0440=>x"AF00",0441=>x"AF00",0442=>x"AF00",0443=>x"AF00",0444=>x"AF00",
0445=>x"AF00",0446=>x"AF00",0447=>x"AF00",0448=>x"AF00",0449=>x"AF00",
0450=>x"AF00",0451=>x"AF00",0452=>x"AF00",0453=>x"AF00",0454=>x"AF00",
0455=>x"AF00",0456=>x"AF00",0457=>x"AF00",0458=>x"AF00",0459=>x"AF00",
0460=>x"AF00",0461=>x"AF00",0462=>x"AF00",0463=>x"AF00",0464=>x"AF00",
0465=>x"AF00",0466=>x"AF00",0467=>x"AF00",0468=>x"AF00",0469=>x"AF00",
0470=>x"AF00",0471=>x"AF00",0472=>x"AF00",0473=>x"AF00",0474=>x"AF00",
0475=>x"AF00",0476=>x"AF00",0477=>x"AF00",0478=>x"AF00",0479=>x"AF00",
0480=>x"AF00",0481=>x"AF00",0482=>x"AF00",0483=>x"AF00",0484=>x"AF00",
0485=>x"AF00",0486=>x"AF00",0487=>x"AF00",0488=>x"AF00",0489=>x"AF00",
0490=>x"AF00",0491=>x"AF00",0492=>x"AF00",0493=>x"AF00",0494=>x"AF00",
0495=>x"AF00",0496=>x"AF00",0497=>x"AF00",0498=>x"AF00",0499=>x"AF00",
0500=>x"AF00",0501=>x"AF00",0502=>x"AF00",0503=>x"AF00",0504=>x"A006",
0505=>x"4800",0506=>x"19FA",0507=>x"AF00",0508=>x"AF00",0509=>x"AF00",
0510=>x"AF00",0511=>x"AF00",0512=>x"5828",0513=>x"5800",0514=>x"5828",
0515=>x"5810",0516=>x"AF00",0517=>x"AF00",0518=>x"AF00",0519=>x"AF00",
0520=>x"AF00",0521=>x"AF00",0522=>x"AF00",0523=>x"AF00",0524=>x"AF00",
0525=>x"AF00",0526=>x"AF00",0527=>x"AF00",0528=>x"AF00",0529=>x"AF00",
0530=>x"AF00",0531=>x"AF00",0532=>x"AF00",0533=>x"AF00",0534=>x"AF00",
0535=>x"AF00",0536=>x"AF00",0537=>x"AF00",0538=>x"AF00",0539=>x"AF00",
0540=>x"AF00",0541=>x"AF00",0542=>x"AF00",0543=>x"AF00",0544=>x"AF00",
0545=>x"AF00",0546=>x"AF00",0547=>x"AF00",0548=>x"AF00",0549=>x"AF00",
0550=>x"AF00",0551=>x"AF00",0552=>x"AF00",0553=>x"AF00",0554=>x"AF00",
0555=>x"AF00",0556=>x"AF00",0557=>x"AF00",0558=>x"AF00",0559=>x"AF00",
0560=>x"AF00",0561=>x"AF00",0562=>x"AF00",0563=>x"AF00",0564=>x"AF00",
0565=>x"AF00",0566=>x"AF00",0567=>x"AF00",0568=>x"AF00",0569=>x"AF00",
0570=>x"AF00",0571=>x"AF00",0572=>x"AF00",0573=>x"AF00",0574=>x"AF00",
0575=>x"AF00",0576=>x"AF00",0577=>x"AF00",0578=>x"AF00",0579=>x"AF00",
0580=>x"AF00",0581=>x"AF00",0582=>x"AF00",0583=>x"AF00",0584=>x"AF00",
0585=>x"AF00",0586=>x"AF00",0587=>x"AF00",0588=>x"AF00",0589=>x"AF00",
0590=>x"AF00",0591=>x"AF00",0592=>x"AF00",0593=>x"AF00",0594=>x"AF00",
0595=>x"AF00",0596=>x"AF00",0597=>x"AF00",0598=>x"AF00",0599=>x"AF00",
0600=>x"AF00",0601=>x"AF00",0602=>x"AF00",0603=>x"AF00",0604=>x"AF00",
0605=>x"AF00",0606=>x"AF00",0607=>x"AF00",0608=>x"AF00",0609=>x"AF00",
0610=>x"AF00",0611=>x"AF00",0612=>x"AF00",0613=>x"AF00",0614=>x"AF00",
0615=>x"AF00",0616=>x"AF00",0617=>x"AF00",0618=>x"AF00",0619=>x"AF00",
0620=>x"AF00",0621=>x"AF00",0622=>x"AF00",0623=>x"AF00",0624=>x"AF00",
0625=>x"AF00",0626=>x"AF00",0627=>x"AF00",0628=>x"AF00",0629=>x"AF00",
0630=>x"AF00",0631=>x"AF00",0632=>x"AF00",0633=>x"AF00",0634=>x"AF00",
0635=>x"AF00",0636=>x"AF00",0637=>x"AF00",0638=>x"AF00",0639=>x"AF00",
0640=>x"AF00",0641=>x"AF00",0642=>x"AF00",0643=>x"AF00",0644=>x"AF00",
0645=>x"AF00",0646=>x"AF00",0647=>x"AF00",0648=>x"AF00",0649=>x"AF00",
0650=>x"AF00",0651=>x"AF00",0652=>x"AF00",0653=>x"AF00",0654=>x"AF00",
0655=>x"AF00",0656=>x"AF00",0657=>x"AF00",0658=>x"AF00",0659=>x"AF00",
0660=>x"AF00",0661=>x"AF00",0662=>x"AF00",0663=>x"AF00",0664=>x"AF00",
0665=>x"AF00",0666=>x"AF00",0667=>x"AF00",0668=>x"AF00",0669=>x"AF00",
0670=>x"AF00",0671=>x"AF00",0672=>x"AF00",0673=>x"AF00",0674=>x"AF00",
0675=>x"AF00",0676=>x"AF00",0677=>x"AF00",0678=>x"AF00",0679=>x"AF00",
0680=>x"AF00",0681=>x"AF00",0682=>x"AF00",0683=>x"AF00",0684=>x"AF00",
0685=>x"AF00",0686=>x"AF00",0687=>x"AF00",0688=>x"AF00",0689=>x"AF00",
0690=>x"AF00",0691=>x"AF00",0692=>x"AF00",0693=>x"AF00",0694=>x"AF00",
0695=>x"AF00",0696=>x"AF00",0697=>x"AF00",0698=>x"AF00",0699=>x"AF00",
0700=>x"AF00",0701=>x"AF00",0702=>x"AF00",0703=>x"AF00",0704=>x"AF00",
0705=>x"AF00",0706=>x"AF00",0707=>x"AF00",0708=>x"AF00",0709=>x"AF00",
0710=>x"AF00",0711=>x"AF00",0712=>x"AF00",0713=>x"AF00",0714=>x"AF00",
0715=>x"AF00",0716=>x"AF00",0717=>x"AF00",0718=>x"AF00",0719=>x"AF00",
0720=>x"AF00",0721=>x"AF00",0722=>x"AF00",0723=>x"AF00",0724=>x"AF00",
0725=>x"AF00",0726=>x"AF00",0727=>x"AF00",0728=>x"AF00",0729=>x"AF00",
0730=>x"AF00",0731=>x"AF00",0732=>x"AF00",0733=>x"AF00",0734=>x"AF00",
0735=>x"AF00",0736=>x"AF00",0737=>x"AF00",0738=>x"AF00",0739=>x"AF00",
0740=>x"AF00",0741=>x"AF00",0742=>x"AF00",0743=>x"AF00",0744=>x"AF00",
0745=>x"AF00",0746=>x"AF00",0747=>x"AF00",0748=>x"AF00",0749=>x"AF00",
0750=>x"AF00",0751=>x"AF00",0752=>x"AF00",0753=>x"AF00",0754=>x"AF00",
0755=>x"AF00",0756=>x"AF00",0757=>x"AF00",0758=>x"AF00",0759=>x"AF00",
0760=>x"A008",0761=>x"4800",0762=>x"19FA",0763=>x"AF00",0764=>x"AF00",
0765=>x"AF00",0766=>x"AF00",0767=>x"AF00",0768=>x"5828",0769=>x"5908",
0770=>x"AF00",0771=>x"AF00",0772=>x"AF00",0773=>x"AF00",0774=>x"AF00",
0775=>x"AF00",0776=>x"AF00",0777=>x"AF00",0778=>x"AF00",0779=>x"AF00",
0780=>x"AF00",0781=>x"AF00",0782=>x"AF00",0783=>x"AF00",0784=>x"AF00",
0785=>x"AF00",0786=>x"AF00",0787=>x"AF00",0788=>x"AF00",0789=>x"AF00",
0790=>x"AF00",0791=>x"AF00",0792=>x"AF00",0793=>x"AF00",0794=>x"AF00",
0795=>x"AF00",0796=>x"AF00",0797=>x"AF00",0798=>x"AF00",0799=>x"AF00",
0800=>x"AF00",0801=>x"AF00",0802=>x"AF00",0803=>x"AF00",0804=>x"AF00",
0805=>x"AF00",0806=>x"AF00",0807=>x"AF00",0808=>x"AF00",0809=>x"AF00",
0810=>x"AF00",0811=>x"AF00",0812=>x"AF00",0813=>x"AF00",0814=>x"AF00",
0815=>x"AF00",0816=>x"AF00",0817=>x"AF00",0818=>x"AF00",0819=>x"AF00",
0820=>x"AF00",0821=>x"AF00",0822=>x"AF00",0823=>x"AF00",0824=>x"AF00",
0825=>x"AF00",0826=>x"AF00",0827=>x"AF00",0828=>x"AF00",0829=>x"AF00",
0830=>x"AF00",0831=>x"AF00",0832=>x"AF00",0833=>x"AF00",0834=>x"AF00",
0835=>x"AF00",0836=>x"AF00",0837=>x"AF00",0838=>x"AF00",0839=>x"AF00",
0840=>x"AF00",0841=>x"AF00",0842=>x"AF00",0843=>x"AF00",0844=>x"AF00",
0845=>x"AF00",0846=>x"AF00",0847=>x"AF00",0848=>x"AF00",0849=>x"AF00",
0850=>x"AF00",0851=>x"AF00",0852=>x"AF00",0853=>x"AF00",0854=>x"AF00",
0855=>x"AF00",0856=>x"AF00",0857=>x"AF00",0858=>x"AF00",0859=>x"AF00",
0860=>x"AF00",0861=>x"AF00",0862=>x"AF00",0863=>x"AF00",0864=>x"AF00",
0865=>x"AF00",0866=>x"AF00",0867=>x"AF00",0868=>x"AF00",0869=>x"AF00",
0870=>x"AF00",0871=>x"AF00",0872=>x"AF00",0873=>x"AF00",0874=>x"AF00",
0875=>x"AF00",0876=>x"AF00",0877=>x"AF00",0878=>x"AF00",0879=>x"AF00",
0880=>x"AF00",0881=>x"AF00",0882=>x"AF00",0883=>x"AF00",0884=>x"AF00",
0885=>x"AF00",0886=>x"AF00",0887=>x"AF00",0888=>x"AF00",0889=>x"AF00",
0890=>x"AF00",0891=>x"AF00",0892=>x"AF00",0893=>x"AF00",0894=>x"AF00",
0895=>x"AF00",0896=>x"AF00",0897=>x"AF00",0898=>x"AF00",0899=>x"AF00",
0900=>x"AF00",0901=>x"AF00",0902=>x"AF00",0903=>x"AF00",0904=>x"AF00",
0905=>x"AF00",0906=>x"AF00",0907=>x"AF00",0908=>x"AF00",0909=>x"AF00",
0910=>x"AF00",0911=>x"AF00",0912=>x"AF00",0913=>x"AF00",0914=>x"AF00",
0915=>x"AF00",0916=>x"AF00",0917=>x"AF00",0918=>x"AF00",0919=>x"AF00",
0920=>x"AF00",0921=>x"AF00",0922=>x"AF00",0923=>x"AF00",0924=>x"AF00",
0925=>x"AF00",0926=>x"AF00",0927=>x"AF00",0928=>x"AF00",0929=>x"AF00",
0930=>x"AF00",0931=>x"AF00",0932=>x"AF00",0933=>x"AF00",0934=>x"AF00",
0935=>x"AF00",0936=>x"AF00",0937=>x"AF00",0938=>x"AF00",0939=>x"AF00",
0940=>x"AF00",0941=>x"AF00",0942=>x"AF00",0943=>x"AF00",0944=>x"AF00",
0945=>x"AF00",0946=>x"AF00",0947=>x"AF00",0948=>x"AF00",0949=>x"AF00",
0950=>x"AF00",0951=>x"AF00",0952=>x"AF00",0953=>x"AF00",0954=>x"AF00",
0955=>x"AF00",0956=>x"AF00",0957=>x"AF00",0958=>x"AF00",0959=>x"AF00",
0960=>x"AF00",0961=>x"AF00",0962=>x"AF00",0963=>x"AF00",0964=>x"AF00",
0965=>x"AF00",0966=>x"AF00",0967=>x"AF00",0968=>x"AF00",0969=>x"AF00",
0970=>x"AF00",0971=>x"AF00",0972=>x"AF00",0973=>x"AF00",0974=>x"AF00",
0975=>x"AF00",0976=>x"AF00",0977=>x"AF00",0978=>x"AF00",0979=>x"AF00",
0980=>x"AF00",0981=>x"AF00",0982=>x"AF00",0983=>x"AF00",0984=>x"AF00",
0985=>x"AF00",0986=>x"AF00",0987=>x"AF00",0988=>x"AF00",0989=>x"AF00",
0990=>x"AF00",0991=>x"AF00",0992=>x"AF00",0993=>x"AF00",0994=>x"AF00",
0995=>x"AF00",0996=>x"AF00",0997=>x"AF00",0998=>x"AF00",0999=>x"AF00",
1000=>x"AF00",1001=>x"AF00",1002=>x"AF00",1003=>x"AF00",1004=>x"AF00",
1005=>x"AF00",1006=>x"AF00",1007=>x"AF00",1008=>x"AF00",1009=>x"AF00",
1010=>x"AF00",1011=>x"AF00",1012=>x"AF00",1013=>x"AF00",1014=>x"AF00",
1015=>x"AF00",1016=>x"A00A",1017=>x"4800",1018=>x"195A",1019=>x"AF00",
1020=>x"AF00",1021=>x"AF00",1022=>x"AF00",1023=>x"AF00",1024=>x"6F01",
1025=>x"5822",1026=>x"6006",1027=>x"C002",1028=>x"5822",1029=>x"6806",
1030=>x"6701",1031=>x"0900",1032=>x"6F01",1033=>x"6F23",1034=>x"0E18",
1035=>x"F816",1036=>x"0034",1037=>x"5F21",1038=>x"E000",1039=>x"C220",
1040=>x"010D",1041=>x"6701",1042=>x"6723",1043=>x"0900",1044=>x"A020",
1045=>x"0F20",1046=>x"0F20",1047=>x"A122",1048=>x"0F3F",1049=>x"5822",
1050=>x"6020",1051=>x"0154",1052=>x"5822",1053=>x"C040",1054=>x"020D",
1055=>x"C022",1056=>x"5822",1057=>x"6820",1058=>x"582E",1059=>x"5D13",
1060=>x"AF00",1061=>x"AF00",1062=>x"AF00",1063=>x"AF00",1064=>x"AF00",
1065=>x"AF00",1066=>x"AF00",1067=>x"AF00",1068=>x"AF00",1069=>x"AF00",
1070=>x"AF00",1071=>x"AF00",1072=>x"AF00",1073=>x"AF00",1074=>x"AF00",
1075=>x"AF00",1076=>x"AF00",1077=>x"AF00",1078=>x"AF00",1079=>x"AF00",
1080=>x"AF00",1081=>x"AF00",1082=>x"AF00",1083=>x"AF00",1084=>x"AF00",
1085=>x"AF00",1086=>x"AF00",1087=>x"AF00",1088=>x"AF00",1089=>x"AF00",
1090=>x"AF00",1091=>x"AF00",1092=>x"AF00",1093=>x"AF00",1094=>x"AF00",
1095=>x"AF00",1096=>x"AF00",1097=>x"AF00",1098=>x"AF00",1099=>x"AF00",
1100=>x"AF00",1101=>x"AF00",1102=>x"AF00",1103=>x"AF00",1104=>x"AF00",
1105=>x"AF00",1106=>x"AF00",1107=>x"AF00",1108=>x"AF00",1109=>x"AF00",
1110=>x"AF00",1111=>x"AF00",1112=>x"AF00",1113=>x"AF00",1114=>x"AF00",
1115=>x"AF00",1116=>x"AF00",1117=>x"AF00",1118=>x"AF00",1119=>x"AF00",
1120=>x"AF00",1121=>x"AF00",1122=>x"AF00",1123=>x"AF00",1124=>x"AF00",
1125=>x"AF00",1126=>x"AF00",1127=>x"AF00",1128=>x"AF00",1129=>x"AF00",
1130=>x"AF00",1131=>x"AF00",1132=>x"AF00",1133=>x"AF00",1134=>x"AF00",
1135=>x"AF00",1136=>x"AF00",1137=>x"AF00",1138=>x"AF00",1139=>x"AF00",
1140=>x"AF00",1141=>x"AF00",1142=>x"AF00",1143=>x"AF00",1144=>x"AF00",
1145=>x"AF00",1146=>x"AF00",1147=>x"AF00",1148=>x"AF00",1149=>x"AF00",
1150=>x"AF00",1151=>x"AF00",1152=>x"AF00",1153=>x"AF00",1154=>x"AF00",
1155=>x"AF00",1156=>x"AF00",1157=>x"AF00",1158=>x"AF00",1159=>x"AF00",
1160=>x"AF00",1161=>x"AF00",1162=>x"AF00",1163=>x"AF00",1164=>x"AF00",
1165=>x"AF00",1166=>x"AF00",1167=>x"AF00",1168=>x"AF00",1169=>x"AF00",
1170=>x"AF00",1171=>x"AF00",1172=>x"AF00",1173=>x"AF00",1174=>x"AF00",
1175=>x"AF00",1176=>x"AF00",1177=>x"AF00",1178=>x"AF00",1179=>x"AF00",
1180=>x"AF00",1181=>x"AF00",1182=>x"AF00",1183=>x"AF00",1184=>x"AF00",
1185=>x"AF00",1186=>x"AF00",1187=>x"AF00",1188=>x"AF00",1189=>x"AF00",
1190=>x"AF00",1191=>x"AF00",1192=>x"A00C",1193=>x"4800",1194=>x"18AA",
1195=>x"AF00",1196=>x"AF00",1197=>x"AF00",1198=>x"AF00",1199=>x"AF00",
1200=>x"AF00",1201=>x"AF00",1202=>x"AF00",1203=>x"AF00",1204=>x"AF00",
1205=>x"AF00",1206=>x"AF00",1207=>x"AF00",1208=>x"AF00",1209=>x"AF00",
1210=>x"AF00",1211=>x"AF00",1212=>x"AF00",1213=>x"AF00",1214=>x"AF00",
1215=>x"AF00",1216=>x"AF00",1217=>x"AF00",1218=>x"AF00",1219=>x"AF00",
1220=>x"AF00",1221=>x"AF00",1222=>x"AF00",1223=>x"AF00",1224=>x"AF00",
1225=>x"AF00",1226=>x"AF00",1227=>x"AF00",1228=>x"AF00",1229=>x"AF00",
1230=>x"AF00",1231=>x"AF00",1232=>x"AF00",1233=>x"AF00",1234=>x"AF00",
1235=>x"AF00",1236=>x"AF00",1237=>x"AF00",1238=>x"AF00",1239=>x"AF00",
1240=>x"AF00",1241=>x"AF00",1242=>x"AF00",1243=>x"AF00",1244=>x"AF00",
1245=>x"AF00",1246=>x"AF00",1247=>x"AF00",1248=>x"AF00",1249=>x"AF00",
1250=>x"AF00",1251=>x"AF00",1252=>x"AF00",1253=>x"AF00",1254=>x"AF00",
1255=>x"AF00",1256=>x"AF00",1257=>x"AF00",1258=>x"AF00",1259=>x"AF00",
1260=>x"AF00",1261=>x"AF00",1262=>x"AF00",1263=>x"AF00",1264=>x"AF00",
1265=>x"AF00",1266=>x"AF00",1267=>x"AF00",1268=>x"AF00",1269=>x"AF00",
1270=>x"AF00",1271=>x"AF00",1272=>x"AF00",1273=>x"AF00",1274=>x"AF00",
1275=>x"AF00",1276=>x"AF00",1277=>x"AF00",1278=>x"AF00",1279=>x"AF00",
1280=>x"A01E",1281=>x"4800",1282=>x"19FA",1283=>x"AF00",1284=>x"AF00",
1285=>x"AF00",1286=>x"AF00",1287=>x"AF00",1288=>x"AF00",1289=>x"AF00",
1290=>x"AF00",1291=>x"AF00",1292=>x"AF00",1293=>x"AF00",1294=>x"AF00",
1295=>x"AF00",1296=>x"AF00",1297=>x"AF00",1298=>x"AF00",1299=>x"AF00",
1300=>x"AF00",1301=>x"AF00",1302=>x"AF00",1303=>x"AF00",1304=>x"AF00",
1305=>x"AF00",1306=>x"AF00",1307=>x"AF00",1308=>x"AF00",1309=>x"AF00",
1310=>x"AF00",1311=>x"AF00",1312=>x"AF00",1313=>x"AF00",1314=>x"AF00",
1315=>x"AF00",1316=>x"AF00",1317=>x"AF00",1318=>x"AF00",1319=>x"AF00",
1320=>x"AF00",1321=>x"AF00",1322=>x"AF00",1323=>x"AF00",1324=>x"AF00",
1325=>x"AF00",1326=>x"AF00",1327=>x"AF00",1328=>x"AF00",1329=>x"AF00",
1330=>x"AF00",1331=>x"AF00",1332=>x"AF00",1333=>x"AF00",1334=>x"AF00",
1335=>x"AF00",1336=>x"AF00",1337=>x"AF00",1338=>x"AF00",1339=>x"AF00",
1340=>x"AF00",1341=>x"AF00",1342=>x"AF00",1343=>x"AF00",1344=>x"AF00",
1345=>x"AF00",1346=>x"AF00",1347=>x"AF00",1348=>x"AF00",1349=>x"AF00",
1350=>x"AF00",1351=>x"AF00",1352=>x"AF00",1353=>x"AF00",1354=>x"AF00",
1355=>x"AF00",1356=>x"AF00",1357=>x"AF00",1358=>x"AF00",1359=>x"AF00",
1360=>x"AF00",1361=>x"AF00",1362=>x"AF00",1363=>x"AF00",1364=>x"AF00",
1365=>x"AF00",1366=>x"AF00",1367=>x"AF00",1368=>x"AF00",1369=>x"AF00",
1370=>x"AF00",1371=>x"AF00",1372=>x"AF00",1373=>x"AF00",1374=>x"AF00",
1375=>x"AF00",1376=>x"AF00",1377=>x"AF00",1378=>x"AF00",1379=>x"AF00",
1380=>x"AF00",1381=>x"AF00",1382=>x"AF00",1383=>x"AF00",1384=>x"AF00",
1385=>x"AF00",1386=>x"AF00",1387=>x"AF00",1388=>x"AF00",1389=>x"AF00",
1390=>x"AF00",1391=>x"AF00",1392=>x"AF00",1393=>x"AF00",1394=>x"AF00",
1395=>x"AF00",1396=>x"AF00",1397=>x"AF00",1398=>x"AF00",1399=>x"AF00",
1400=>x"AF00",1401=>x"AF00",1402=>x"AF00",1403=>x"AF00",1404=>x"AF00",
1405=>x"AF00",1406=>x"AF00",1407=>x"AF00",1408=>x"AF00",1409=>x"AF00",
1410=>x"AF00",1411=>x"AF00",1412=>x"AF00",1413=>x"AF00",1414=>x"AF00",
1415=>x"AF00",1416=>x"AF00",1417=>x"AF00",1418=>x"AF00",1419=>x"AF00",
1420=>x"AF00",1421=>x"AF00",1422=>x"AF00",1423=>x"AF00",1424=>x"AF00",
1425=>x"AF00",1426=>x"AF00",1427=>x"AF00",1428=>x"AF00",1429=>x"AF00",
1430=>x"AF00",1431=>x"AF00",1432=>x"AF00",1433=>x"AF00",1434=>x"AF00",
1435=>x"AF00",1436=>x"AF00",1437=>x"AF00",1438=>x"AF00",1439=>x"AF00",
1440=>x"AF00",1441=>x"AF00",1442=>x"AF00",1443=>x"AF00",1444=>x"AF00",
1445=>x"AF00",1446=>x"AF00",1447=>x"AF00",1448=>x"AF00",1449=>x"AF00",
1450=>x"AF00",1451=>x"AF00",1452=>x"AF00",1453=>x"AF00",1454=>x"AF00",
1455=>x"AF00",1456=>x"AF00",1457=>x"AF00",1458=>x"AF00",1459=>x"AF00",
1460=>x"AF00",1461=>x"AF00",1462=>x"AF00",1463=>x"AF00",1464=>x"AF00",
1465=>x"AF00",1466=>x"AF00",1467=>x"AF00",1468=>x"AF00",1469=>x"AF00",
1470=>x"AF00",1471=>x"AF00",1472=>x"AF00",1473=>x"AF00",1474=>x"AF00",
1475=>x"AF00",1476=>x"AF00",1477=>x"AF00",1478=>x"AF00",1479=>x"AF00",
1480=>x"AF00",1481=>x"AF00",1482=>x"AF00",1483=>x"AF00",1484=>x"AF00",
1485=>x"AF00",1486=>x"AF00",1487=>x"AF00",1488=>x"AF00",1489=>x"AF00",
1490=>x"AF00",1491=>x"AF00",1492=>x"AF00",1493=>x"AF00",1494=>x"AF00",
1495=>x"AF00",1496=>x"AF00",1497=>x"AF00",1498=>x"AF00",1499=>x"AF00",
1500=>x"AF00",1501=>x"AF00",1502=>x"AF00",1503=>x"AF00",1504=>x"AF00",
1505=>x"AF00",1506=>x"AF00",1507=>x"AF00",1508=>x"AF00",1509=>x"AF00",
1510=>x"AF00",1511=>x"AF00",1512=>x"AF00",1513=>x"AF00",1514=>x"AF00",
1515=>x"AF00",1516=>x"AF00",1517=>x"AF00",1518=>x"AF00",1519=>x"AF00",
1520=>x"AF00",1521=>x"AF00",1522=>x"AF00",1523=>x"AF00",1524=>x"AF00",
1525=>x"AF00",1526=>x"AF00",1527=>x"AF00",1528=>x"AF00",1529=>x"AF00",
1530=>x"AF00",1531=>x"AF00",1532=>x"AF00",1533=>x"AF00",1534=>x"AF00",
1535=>x"AF00",1536=>x"A010",1537=>x"4800",1538=>x"19AA",1539=>x"AF00",
1540=>x"AF00",1541=>x"AF00",1542=>x"AF00",1543=>x"AF00",1544=>x"AF00",
1545=>x"AF00",1546=>x"AF00",1547=>x"AF00",1548=>x"AF00",1549=>x"AF00",
1550=>x"AF00",1551=>x"AF00",1552=>x"AF00",1553=>x"AF00",1554=>x"AF00",
1555=>x"AF00",1556=>x"AF00",1557=>x"AF00",1558=>x"AF00",1559=>x"AF00",
1560=>x"AF00",1561=>x"AF00",1562=>x"AF00",1563=>x"AF00",1564=>x"AF00",
1565=>x"AF00",1566=>x"AF00",1567=>x"AF00",1568=>x"AF00",1569=>x"AF00",
1570=>x"AF00",1571=>x"AF00",1572=>x"AF00",1573=>x"AF00",1574=>x"AF00",
1575=>x"AF00",1576=>x"AF00",1577=>x"AF00",1578=>x"AF00",1579=>x"AF00",
1580=>x"AF00",1581=>x"AF00",1582=>x"AF00",1583=>x"AF00",1584=>x"AF00",
1585=>x"AF00",1586=>x"AF00",1587=>x"AF00",1588=>x"AF00",1589=>x"AF00",
1590=>x"AF00",1591=>x"AF00",1592=>x"AF00",1593=>x"AF00",1594=>x"AF00",
1595=>x"AF00",1596=>x"AF00",1597=>x"AF00",1598=>x"AF00",1599=>x"AF00",
1600=>x"AF00",1601=>x"AF00",1602=>x"AF00",1603=>x"AF00",1604=>x"AF00",
1605=>x"AF00",1606=>x"AF00",1607=>x"AF00",1608=>x"AF00",1609=>x"AF00",
1610=>x"AF00",1611=>x"AF00",1612=>x"AF00",1613=>x"AF00",1614=>x"AF00",
1615=>x"AF00",1616=>x"AF00",1617=>x"AF00",1618=>x"AF00",1619=>x"AF00",
1620=>x"AF00",1621=>x"AF00",1622=>x"AF00",1623=>x"AF00",1624=>x"AF00",
1625=>x"AF00",1626=>x"AF00",1627=>x"AF00",1628=>x"AF00",1629=>x"AF00",
1630=>x"AF00",1631=>x"AF00",1632=>x"AF00",1633=>x"AF00",1634=>x"AF00",
1635=>x"AF00",1636=>x"AF00",1637=>x"AF00",1638=>x"AF00",1639=>x"AF00",
1640=>x"AF00",1641=>x"AF00",1642=>x"AF00",1643=>x"AF00",1644=>x"AF00",
1645=>x"AF00",1646=>x"AF00",1647=>x"AF00",1648=>x"AF00",1649=>x"AF00",
1650=>x"AF00",1651=>x"AF00",1652=>x"AF00",1653=>x"AF00",1654=>x"AF00",
1655=>x"AF00",1656=>x"AF00",1657=>x"AF00",1658=>x"AF00",1659=>x"AF00",
1660=>x"AF00",1661=>x"AF00",1662=>x"AF00",1663=>x"AF00",1664=>x"AF00",
1665=>x"AF00",1666=>x"AF00",1667=>x"AF00",1668=>x"AF00",1669=>x"AF00",
1670=>x"AF00",1671=>x"AF00",1672=>x"AF00",1673=>x"AF00",1674=>x"AF00",
1675=>x"AF00",1676=>x"AF00",1677=>x"AF00",1678=>x"AF00",1679=>x"AF00",
1680=>x"AF00",1681=>x"AF00",1682=>x"AF00",1683=>x"AF00",1684=>x"AF00",
1685=>x"AF00",1686=>x"AF00",1687=>x"AF00",1688=>x"AF00",1689=>x"AF00",
1690=>x"AF00",1691=>x"AF00",1692=>x"AF00",1693=>x"AF00",1694=>x"AF00",
1695=>x"AF00",1696=>x"AF00",1697=>x"AF00",1698=>x"AF00",1699=>x"AF00",
1700=>x"AF00",1701=>x"AF00",1702=>x"AF00",1703=>x"AF00",1704=>x"AF00",
1705=>x"AF00",1706=>x"AF00",1707=>x"AF00",1708=>x"AF00",1709=>x"AF00",
1710=>x"AF00",1711=>x"AF00",1712=>x"AF00",1713=>x"AF00",1714=>x"AF00",
1715=>x"AF00",1716=>x"AF00",1717=>x"AF00",1718=>x"AF00",1719=>x"AF00",
1720=>x"AF00",1721=>x"AF00",1722=>x"AF00",1723=>x"AF00",1724=>x"AF00",
1725=>x"AF00",1726=>x"AF00",1727=>x"AF00",1728=>x"AF00",1729=>x"AF00",
1730=>x"AF00",1731=>x"AF00",1732=>x"AF00",1733=>x"AF00",1734=>x"AF00",
1735=>x"AF00",1736=>x"AF00",1737=>x"AF00",1738=>x"AF00",1739=>x"AF00",
1740=>x"AF00",1741=>x"AF00",1742=>x"AF00",1743=>x"AF00",1744=>x"AF00",
1745=>x"AF00",1746=>x"AF00",1747=>x"AF00",1748=>x"AF00",1749=>x"AF00",
1750=>x"AF00",1751=>x"AF00",1752=>x"A012",1753=>x"4800",1754=>x"183A",
1755=>x"AF00",1756=>x"AF00",1757=>x"AF00",1758=>x"AF00",1759=>x"AF00",
1760=>x"5820",1761=>x"A0FE",1762=>x"C8E2",1763=>x"2FE3",1764=>x"AF00",
1765=>x"AC00",1766=>x"02AA",1767=>x"17F1",1768=>x"4824",1769=>x"17ED",
1770=>x"4802",1771=>x"17E9",1772=>x"A042",1773=>x"4846",1774=>x"17E3",
1775=>x"A040",1776=>x"4846",1777=>x"17DD",1778=>x"054B",1779=>x"A2F4",
1780=>x"48E0",1781=>x"AC00",1782=>x"AF00",1783=>x"AF00",1784=>x"A014",
1785=>x"4800",1786=>x"19BC",1787=>x"AF00",1788=>x"AF00",1789=>x"A2FE",
1790=>x"48E0",1791=>x"AF00",1792=>x"A000",1793=>x"A0C0",1794=>x"4804",
1795=>x"4806",1796=>x"A310",1797=>x"A020",1798=>x"17BF",1799=>x"A648",
1800=>x"17AF",1801=>x"C842",1802=>x"2FD3",1803=>x"A062",1804=>x"A310",
1805=>x"17B1",1806=>x"A054",1807=>x"17A1",1808=>x"C842",1809=>x"2FD3",
1810=>x"C862",1811=>x"2F87",1812=>x"A018",1813=>x"17A1",1814=>x"A002",
1815=>x"179D",1816=>x"A00C",1817=>x"1799",1818=>x"A022",1819=>x"AF00",
1820=>x"A500",1821=>x"1791",1822=>x"A504",1823=>x"178D",1824=>x"A41E",
1825=>x"1789",1826=>x"A40E",1827=>x"1785",1828=>x"A200",1829=>x"1781",
1830=>x"A300",1831=>x"177D",1832=>x"A314",1833=>x"1779",1834=>x"A200",
1835=>x"1775",1836=>x"5822",1837=>x"6042",1838=>x"8854",1839=>x"2868",
1840=>x"0214",1841=>x"C814",1842=>x"C854",1843=>x"C300",1844=>x"1763",
1845=>x"1804",1846=>x"A200",1847=>x"175D",1848=>x"0214",1849=>x"C300",
1850=>x"1757",1851=>x"A020",1852=>x"A401",1853=>x"1751",1854=>x"AF00",
1855=>x"A022",1856=>x"A500",1857=>x"1749",1858=>x"A504",1859=>x"1745",
1860=>x"AF00",1861=>x"AF00",1862=>x"AF00",1863=>x"AF00",1864=>x"A41E",
1865=>x"1739",1866=>x"A40E",1867=>x"1735",1868=>x"A200",1869=>x"1731",
1870=>x"A302",1871=>x"172D",1872=>x"A314",1873=>x"1729",1874=>x"A200",
1875=>x"1725",1876=>x"5822",1877=>x"6044",1878=>x"8854",1879=>x"2868",
1880=>x"0214",1881=>x"C814",1882=>x"C854",1883=>x"C300",1884=>x"1713",
1885=>x"1804",1886=>x"A200",1887=>x"170D",1888=>x"0214",1889=>x"C300",
1890=>x"1707",1891=>x"1820",1892=>x"AF00",1893=>x"AF00",1894=>x"AF00",
1895=>x"AF00",1896=>x"AF00",1897=>x"AF00",1898=>x"AF00",1899=>x"AF00",
1900=>x"AF00",1901=>x"AF00",1902=>x"AF00",1903=>x"AF00",1904=>x"AF00",
1905=>x"AF00",1906=>x"AF00",1907=>x"AF00",1908=>x"A2FA",1909=>x"48E0",
1910=>x"0B00",1911=>x"1FFF",1912=>x"AF00",1913=>x"AF00",1914=>x"AF00",
1915=>x"AF00",1916=>x"AF00",1917=>x"AF00",1918=>x"AF00",1919=>x"AF00",
1920=>x"AF00",1921=>x"AF00",1922=>x"AF00",1923=>x"AF00",1924=>x"AF00",
1925=>x"AF00",1926=>x"AF00",1927=>x"AF00",1928=>x"AF00",1929=>x"AF00",
1930=>x"AF00",1931=>x"AF00",1932=>x"AF00",1933=>x"AF00",1934=>x"AF00",
1935=>x"AF00",1936=>x"AF00",1937=>x"AF00",1938=>x"AF00",1939=>x"AF00",
1940=>x"AF00",1941=>x"AF00",1942=>x"AF00",1943=>x"AF00",1944=>x"AF00",
1945=>x"AF00",1946=>x"AF00",1947=>x"AF00",1948=>x"AF00",1949=>x"AF00",
1950=>x"AF00",1951=>x"AF00",1952=>x"AF00",1953=>x"AF00",1954=>x"AF00",
1955=>x"AF00",1956=>x"AF00",1957=>x"AF00",1958=>x"AF00",1959=>x"AF00",
1960=>x"AF00",1961=>x"AF00",1962=>x"AF00",1963=>x"AF00",1964=>x"AF00",
1965=>x"AF00",1966=>x"AF00",1967=>x"AF00",1968=>x"AF00",1969=>x"AF00",
1970=>x"AF00",1971=>x"AF00",1972=>x"AF00",1973=>x"AF00",1974=>x"AF00",
1975=>x"AF00",1976=>x"AF00",1977=>x"AF00",1978=>x"AF00",1979=>x"AF00",
1980=>x"AF00",1981=>x"AF00",1982=>x"AF00",1983=>x"AF00",1984=>x"AF00",
1985=>x"AF00",1986=>x"AF00",1987=>x"AF00",1988=>x"AF00",1989=>x"AF00",
1990=>x"AF00",1991=>x"AF00",1992=>x"AF00",1993=>x"AF00",1994=>x"AF00",
1995=>x"AF00",1996=>x"AF00",1997=>x"AF00",1998=>x"AF00",1999=>x"AF00",
2000=>x"AF00",2001=>x"AF00",2002=>x"AF00",2003=>x"AF00",2004=>x"AF00",
2005=>x"AF00",2006=>x"AF00",2007=>x"AF00",2008=>x"AF00",2009=>x"A000",
2010=>x"4800",2011=>x"AF00",2012=>x"5822",2013=>x"6000",2014=>x"0F00",
2015=>x"A120",2016=>x"A042",2017=>x"8804",2018=>x"2894",2019=>x"8806",
2020=>x"28F4",2021=>x"5F21",2022=>x"A002",2023=>x"6A02",2024=>x"0F3F",
2025=>x"0F5F",2026=>x"5830",2027=>x"5800",2028=>x"5F21",2029=>x"A004",
2030=>x"6A02",2031=>x"0F3F",2032=>x"0F5F",2033=>x"5830",2034=>x"5800",
2035=>x"AF00",2036=>x"5822",2037=>x"6002",2038=>x"5822",2039=>x"6024",
2040=>x"1E09",2041=>x"AF00",2042=>x"AF00",2043=>x"AF00",2044=>x"A008",
2045=>x"0F1F",2046=>x"A000",2047=>x"A022",2048=>x"A0EE",2049=>x"88E0",
2050=>x"286C",2051=>x"AF00",2052=>x"0054",2053=>x"0114",2054=>x"0238",
2055=>x"C8E2",2056=>x"2FB7",2057=>x"AF00",2058=>x"A0F4",2059=>x"48E0",
2060=>x"0801",2061=>x"AF00",2062=>x"AF00",2063=>x"AF00",2064=>x"AF00",
2065=>x"AF00",2066=>x"AF00",2067=>x"AF00",2068=>x"AF00",2069=>x"AF00",
2070=>x"AF00",2071=>x"AF00",2072=>x"AF00",2073=>x"AF00",2074=>x"AF00",
2075=>x"AF00",2076=>x"AF00",2077=>x"AF00",2078=>x"AF00",2079=>x"AF00",
2080=>x"AF00",2081=>x"AF00",2082=>x"AF00",2083=>x"AF00",2084=>x"AF00",
2085=>x"AF00",2086=>x"AF00",2087=>x"AF00",2088=>x"AF00",2089=>x"AF00",
2090=>x"AF00",2091=>x"AF00",2092=>x"AF00",2093=>x"AF00",2094=>x"AF00",
2095=>x"AF00",2096=>x"AF00",2097=>x"AF00",2098=>x"AF00",2099=>x"AF00",
2100=>x"AF00",2101=>x"AF00",2102=>x"AF00",2103=>x"AF00",2104=>x"AF00",
2105=>x"AF00",2106=>x"AF00",2107=>x"AF00",2108=>x"AF00",2109=>x"AF00",
2110=>x"AF00",2111=>x"AF00",2112=>x"AF00",2113=>x"AF00",2114=>x"AF00",
2115=>x"AF00",2116=>x"AF00",2117=>x"AF00",2118=>x"AF00",2119=>x"AF00",
2120=>x"AF00",2121=>x"AF00",2122=>x"AF00",2123=>x"AF00",2124=>x"AF00",
2125=>x"AF00",2126=>x"AF00",2127=>x"AF00",2128=>x"AF00",2129=>x"AF00",
2130=>x"AF00",2131=>x"AF00",2132=>x"AF00",2133=>x"AF00",2134=>x"AF00",
2135=>x"AF00",2136=>x"AF00",2137=>x"AF00",2138=>x"AF00",2139=>x"AF00",
2140=>x"AF00",2141=>x"AF00",2142=>x"AF00",2143=>x"AF00",2144=>x"AF00",
2145=>x"AF00",2146=>x"AF00",2147=>x"AF00",2148=>x"AF00",2149=>x"AF00",
2150=>x"AF00",2151=>x"AF00",2152=>x"AF00",2153=>x"AF00",2154=>x"AF00",
2155=>x"AF00",2156=>x"AF00",2157=>x"AF00",2158=>x"AF00",2159=>x"AF00",
2160=>x"AF00",2161=>x"AF00",2162=>x"AF00",2163=>x"AF00",2164=>x"AF00",
2165=>x"AF00",2166=>x"AF00",2167=>x"AF00",2168=>x"AF00",2169=>x"AF00",
2170=>x"AF00",2171=>x"AF00",2172=>x"AF00",2173=>x"AF00",2174=>x"AF00",
2175=>x"AF00",2176=>x"AF00",2177=>x"AF00",2178=>x"AF00",2179=>x"AF00",
2180=>x"AF00",2181=>x"AF00",2182=>x"AF00",2183=>x"AF00",2184=>x"AF00",
2185=>x"AF00",2186=>x"AF00",2187=>x"AF00",2188=>x"AF00",2189=>x"AF00",
2190=>x"AF00",2191=>x"AF00",2192=>x"AF00",2193=>x"AF00",2194=>x"AF00",
2195=>x"AF00",2196=>x"AF00",2197=>x"AF00",2198=>x"AF00",2199=>x"AF00",
2200=>x"AF00",2201=>x"AF00",2202=>x"AF00",2203=>x"AF00",2204=>x"AF00",
2205=>x"AF00",2206=>x"AF00",2207=>x"AF00",2208=>x"AF00",2209=>x"AF00",
2210=>x"AF00",2211=>x"AF00",2212=>x"AF00",2213=>x"AF00",2214=>x"AF00",
2215=>x"AF00",2216=>x"AF00",2217=>x"AF00",2218=>x"AF00",2219=>x"AF00",
2220=>x"AF00",2221=>x"AF00",2222=>x"AF00",2223=>x"AF00",2224=>x"AF00",
2225=>x"AF00",2226=>x"AF00",2227=>x"AF00",2228=>x"AF00",2229=>x"AF00",
2230=>x"AF00",2231=>x"AF00",2232=>x"AF00",2233=>x"AF00",2234=>x"AF00",
2235=>x"AF00",2236=>x"AF00",2237=>x"AF00",2238=>x"AF00",2239=>x"AF00",
2240=>x"AF00",2241=>x"AF00",2242=>x"AF00",2243=>x"AF00",2244=>x"AF00",
2245=>x"AF00",2246=>x"AF00",2247=>x"AF00",2248=>x"AF00",2249=>x"AF00",
2250=>x"AF00",2251=>x"AF00",2252=>x"AF00",2253=>x"AF00",2254=>x"AF00",
2255=>x"AF00",2256=>x"AF00",2257=>x"AF00",2258=>x"AF00",2259=>x"AF00",
2260=>x"AF00",2261=>x"AF00",2262=>x"AF00",2263=>x"AF00",2264=>x"AF00",
2265=>x"AF00",2266=>x"AF00",2267=>x"AF00",2268=>x"AF00",2269=>x"AF00",
2270=>x"AF00",2271=>x"AF00",2272=>x"AF00",2273=>x"AF00",2274=>x"AF00",
2275=>x"AF00",2276=>x"AF00",2277=>x"AF00",2278=>x"AF00",2279=>x"AF00",
2280=>x"AF00",2281=>x"AF00",2282=>x"AF00",2283=>x"AF00",2284=>x"AF00",
2285=>x"AF00",2286=>x"AF00",2287=>x"AF00",2288=>x"AF00",2289=>x"AF00",
2290=>x"AF00",2291=>x"AF00",2292=>x"AF00",2293=>x"AF00",2294=>x"AF00",
2295=>x"AF00",2296=>x"AF00",2297=>x"AF00",2298=>x"AF00",2299=>x"AF00",
2300=>x"AF00",2301=>x"AF00",2302=>x"AF00",2303=>x"AF00",2304=>x"AF00",
2305=>x"AF00",2306=>x"AF00",2307=>x"AF00",2308=>x"AF00",2309=>x"AF00",
2310=>x"AF00",2311=>x"AF00",2312=>x"AF00",2313=>x"AF00",2314=>x"AF00",
2315=>x"AF00",2316=>x"AF00",2317=>x"AF00",2318=>x"AF00",2319=>x"AF00",
2320=>x"AF00",2321=>x"AF00",2322=>x"AF00",2323=>x"AF00",2324=>x"AF00",
2325=>x"AF00",2326=>x"AF00",2327=>x"AF00",2328=>x"AF00",2329=>x"AF00",
2330=>x"AF00",2331=>x"AF00",2332=>x"AF00",2333=>x"AF00",2334=>x"AF00",
2335=>x"AF00",2336=>x"AF00",2337=>x"AF00",2338=>x"AF00",2339=>x"AF00",
2340=>x"AF00",2341=>x"AF00",2342=>x"AF00",2343=>x"AF00",2344=>x"AF00",
2345=>x"AF00",2346=>x"AF00",2347=>x"AF00",2348=>x"AF00",2349=>x"AF00",
2350=>x"AF00",2351=>x"AF00",2352=>x"AF00",2353=>x"AF00",2354=>x"AF00",
2355=>x"AF00",2356=>x"AF00",2357=>x"AF00",2358=>x"AF00",2359=>x"AF00",
2360=>x"AF00",2361=>x"AF00",2362=>x"AF00",2363=>x"AF00",2364=>x"AF00",
2365=>x"AF00",2366=>x"AF00",2367=>x"AF00",2368=>x"AF00",2369=>x"AF00",
2370=>x"AF00",2371=>x"AF00",2372=>x"AF00",2373=>x"AF00",2374=>x"AF00",
2375=>x"AF00",2376=>x"AF00",2377=>x"AF00",2378=>x"AF00",2379=>x"AF00",
2380=>x"AF00",2381=>x"AF00",2382=>x"AF00",2383=>x"AF00",2384=>x"AF00",
2385=>x"AF00",2386=>x"AF00",2387=>x"AF00",2388=>x"AF00",2389=>x"AF00",
2390=>x"AF00",2391=>x"AF00",2392=>x"AF00",2393=>x"AF00",2394=>x"AF00",
2395=>x"AF00",2396=>x"AF00",2397=>x"AF00",2398=>x"AF00",2399=>x"AF00",
2400=>x"AF00",2401=>x"AF00",2402=>x"AF00",2403=>x"AF00",2404=>x"AF00",
2405=>x"AF00",2406=>x"AF00",2407=>x"AF00",2408=>x"AF00",2409=>x"AF00",
2410=>x"AF00",2411=>x"AF00",2412=>x"AF00",2413=>x"AF00",2414=>x"AF00",
2415=>x"AF00",2416=>x"AF00",2417=>x"AF00",2418=>x"AF00",2419=>x"AF00",
2420=>x"AF00",2421=>x"AF00",2422=>x"AF00",2423=>x"AF00",2424=>x"AF00",
2425=>x"AF00",2426=>x"AF00",2427=>x"AF00",2428=>x"AF00",2429=>x"AF00",
2430=>x"AF00",2431=>x"AF00",2432=>x"AF00",2433=>x"AF00",2434=>x"AF00",
2435=>x"AF00",2436=>x"AF00",2437=>x"AF00",2438=>x"AF00",2439=>x"AF00",
2440=>x"AF00",2441=>x"AF00",2442=>x"AF00",2443=>x"AF00",2444=>x"AF00",
2445=>x"AF00",2446=>x"AF00",2447=>x"AF00",2448=>x"AF00",2449=>x"AF00",
2450=>x"AF00",2451=>x"AF00",2452=>x"AF00",2453=>x"AF00",2454=>x"AF00",
2455=>x"AF00",2456=>x"AF00",2457=>x"AF00",2458=>x"AF00",2459=>x"AF00",
2460=>x"AF00",2461=>x"AF00",2462=>x"AF00",2463=>x"AF00",2464=>x"AF00",
2465=>x"AF00",2466=>x"AF00",2467=>x"AF00",2468=>x"AF00",2469=>x"AF00",
2470=>x"AF00",2471=>x"AF00",2472=>x"AF00",2473=>x"AF00",2474=>x"AF00",
2475=>x"AF00",2476=>x"AF00",2477=>x"AF00",2478=>x"AF00",2479=>x"AF00",
2480=>x"AF00",2481=>x"AF00",2482=>x"AF00",2483=>x"AF00",2484=>x"AF00",
2485=>x"AF00",2486=>x"AF00",2487=>x"AF00",2488=>x"AF00",2489=>x"AF00",
2490=>x"AF00",2491=>x"AF00",2492=>x"AF00",2493=>x"AF00",2494=>x"AF00",
2495=>x"AF00",2496=>x"AF00",2497=>x"AF00",2498=>x"AF00",2499=>x"AF00",
2500=>x"AF00",2501=>x"AF00",2502=>x"AF00",2503=>x"AF00",2504=>x"AF00",
2505=>x"AF00",2506=>x"AF00",2507=>x"AF00",2508=>x"AF00",2509=>x"AF00",
2510=>x"AF00",2511=>x"AF00",2512=>x"AF00",2513=>x"AF00",2514=>x"AF00",
2515=>x"AF00",2516=>x"AF00",2517=>x"AF00",2518=>x"AF00",2519=>x"AF00",
2520=>x"AF00",2521=>x"AF00",2522=>x"AF00",2523=>x"AF00",2524=>x"AF00",
2525=>x"AF00",2526=>x"AF00",2527=>x"AF00",2528=>x"AF00",2529=>x"AF00",
2530=>x"AF00",2531=>x"AF00",2532=>x"AF00",2533=>x"AF00",2534=>x"AF00",
2535=>x"AF00",2536=>x"AF00",2537=>x"AF00",2538=>x"AF00",2539=>x"AF00",
2540=>x"AF00",2541=>x"AF00",2542=>x"AF00",2543=>x"AF00",2544=>x"AF00",
2545=>x"AF00",2546=>x"AF00",2547=>x"AF00",2548=>x"AF00",2549=>x"AF00",
2550=>x"AF00",2551=>x"AF00",2552=>x"AF00",2553=>x"AF00",2554=>x"AF00",
2555=>x"AF00",2556=>x"AF00",2557=>x"AF00",2558=>x"AF00",2559=>x"AF00",
2560=>x"AF00",2561=>x"AF00",2562=>x"AF00",2563=>x"AF00",2564=>x"AF00",
2565=>x"AF00",2566=>x"AF00",2567=>x"AF00",2568=>x"AF00",2569=>x"AF00",
2570=>x"AF00",2571=>x"AF00",2572=>x"AF00",2573=>x"AF00",2574=>x"AF00",
2575=>x"AF00",2576=>x"AF00",2577=>x"AF00",2578=>x"AF00",2579=>x"AF00",
2580=>x"AF00",2581=>x"AF00",2582=>x"AF00",2583=>x"AF00",2584=>x"AF00",
2585=>x"AF00",2586=>x"AF00",2587=>x"AF00",2588=>x"AF00",2589=>x"AF00",
2590=>x"AF00",2591=>x"AF00",2592=>x"AF00",2593=>x"AF00",2594=>x"AF00",
2595=>x"AF00",2596=>x"AF00",2597=>x"AF00",2598=>x"AF00",2599=>x"AF00",
2600=>x"AF00",2601=>x"AF00",2602=>x"AF00",2603=>x"AF00",2604=>x"AF00",
2605=>x"AF00",2606=>x"AF00",2607=>x"AF00",2608=>x"AF00",2609=>x"AF00",
2610=>x"AF00",2611=>x"AF00",2612=>x"AF00",2613=>x"AF00",2614=>x"AF00",
2615=>x"AF00",2616=>x"AF00",2617=>x"AF00",2618=>x"AF00",2619=>x"AF00",
2620=>x"AF00",2621=>x"AF00",2622=>x"AF00",2623=>x"AF00",2624=>x"AF00",
2625=>x"AF00",2626=>x"AF00",2627=>x"AF00",2628=>x"AF00",2629=>x"AF00",
2630=>x"AF00",2631=>x"AF00",2632=>x"AF00",2633=>x"AF00",2634=>x"AF00",
2635=>x"AF00",2636=>x"AF00",2637=>x"AF00",2638=>x"AF00",2639=>x"AF00",
2640=>x"AF00",2641=>x"AF00",2642=>x"AF00",2643=>x"AF00",2644=>x"AF00",
2645=>x"AF00",2646=>x"AF00",2647=>x"AF00",2648=>x"AF00",2649=>x"AF00",
2650=>x"AF00",2651=>x"AF00",2652=>x"AF00",2653=>x"AF00",2654=>x"AF00",
2655=>x"AF00",2656=>x"AF00",2657=>x"AF00",2658=>x"AF00",2659=>x"AF00",
2660=>x"AF00",2661=>x"AF00",2662=>x"AF00",2663=>x"AF00",2664=>x"AF00",
2665=>x"AF00",2666=>x"AF00",2667=>x"AF00",2668=>x"AF00",2669=>x"AF00",
2670=>x"AF00",2671=>x"AF00",2672=>x"AF00",2673=>x"AF00",2674=>x"AF00",
2675=>x"AF00",2676=>x"AF00",2677=>x"AF00",2678=>x"AF00",2679=>x"AF00",
2680=>x"AF00",2681=>x"AF00",2682=>x"AF00",2683=>x"AF00",2684=>x"AF00",
2685=>x"AF00",2686=>x"AF00",2687=>x"AF00",2688=>x"AF00",2689=>x"AF00",
2690=>x"AF00",2691=>x"AF00",2692=>x"AF00",2693=>x"AF00",2694=>x"AF00",
2695=>x"AF00",2696=>x"AF00",2697=>x"AF00",2698=>x"AF00",2699=>x"AF00",
2700=>x"AF00",2701=>x"AF00",2702=>x"AF00",2703=>x"AF00",2704=>x"AF00",
2705=>x"AF00",2706=>x"AF00",2707=>x"AF00",2708=>x"AF00",2709=>x"AF00",
2710=>x"AF00",2711=>x"AF00",2712=>x"AF00",2713=>x"AF00",2714=>x"AF00",
2715=>x"AF00",2716=>x"AF00",2717=>x"AF00",2718=>x"AF00",2719=>x"AF00",
2720=>x"AF00",2721=>x"AF00",2722=>x"AF00",2723=>x"AF00",2724=>x"AF00",
2725=>x"AF00",2726=>x"AF00",2727=>x"AF00",2728=>x"AF00",2729=>x"AF00",
2730=>x"AF00",2731=>x"AF00",2732=>x"AF00",2733=>x"AF00",2734=>x"AF00",
2735=>x"AF00",2736=>x"AF00",2737=>x"AF00",2738=>x"AF00",2739=>x"AF00",
2740=>x"AF00",2741=>x"AF00",2742=>x"AF00",2743=>x"AF00",2744=>x"AF00",
2745=>x"AF00",2746=>x"AF00",2747=>x"AF00",2748=>x"AF00",2749=>x"AF00",
2750=>x"AF00",2751=>x"AF00",2752=>x"AF00",2753=>x"AF00",2754=>x"AF00",
2755=>x"AF00",2756=>x"AF00",2757=>x"AF00",2758=>x"AF00",2759=>x"AF00",
2760=>x"AF00",2761=>x"AF00",2762=>x"AF00",2763=>x"AF00",2764=>x"AF00",
2765=>x"AF00",2766=>x"AF00",2767=>x"AF00",2768=>x"AF00",2769=>x"AF00",
2770=>x"AF00",2771=>x"AF00",2772=>x"AF00",2773=>x"AF00",2774=>x"AF00",
2775=>x"AF00",2776=>x"AF00",2777=>x"AF00",2778=>x"AF00",2779=>x"AF00",
2780=>x"AF00",2781=>x"AF00",2782=>x"AF00",2783=>x"AF00",2784=>x"AF00",
2785=>x"AF00",2786=>x"AF00",2787=>x"AF00",2788=>x"AF00",2789=>x"AF00",
2790=>x"AF00",2791=>x"AF00",2792=>x"AF00",2793=>x"AF00",2794=>x"AF00",
2795=>x"AF00",2796=>x"AF00",2797=>x"AF00",2798=>x"AF00",2799=>x"AF00",
2800=>x"AF00",2801=>x"AF00",2802=>x"AF00",2803=>x"AF00",2804=>x"AF00",
2805=>x"AF00",2806=>x"AF00",2807=>x"AF00",2808=>x"AF00",2809=>x"AF00",
2810=>x"AF00",2811=>x"AF00",2812=>x"AF00",2813=>x"AF00",2814=>x"AF00",
2815=>x"AF00",2816=>x"AF00",2817=>x"AF00",2818=>x"AF00",2819=>x"AF00",
2820=>x"AF00",2821=>x"AF00",2822=>x"AF00",2823=>x"AF00",2824=>x"AF00",
2825=>x"AF00",2826=>x"AF00",2827=>x"AF00",2828=>x"AF00",2829=>x"AF00",
2830=>x"AF00",2831=>x"AF00",2832=>x"AF00",2833=>x"AF00",2834=>x"AF00",
2835=>x"AF00",2836=>x"AF00",2837=>x"AF00",2838=>x"AF00",2839=>x"AF00",
2840=>x"AF00",2841=>x"AF00",2842=>x"AF00",2843=>x"AF00",2844=>x"AF00",
2845=>x"AF00",2846=>x"AF00",2847=>x"AF00",2848=>x"AF00",2849=>x"AF00",
2850=>x"AF00",2851=>x"AF00",2852=>x"AF00",2853=>x"AF00",2854=>x"AF00",
2855=>x"AF00",2856=>x"AF00",2857=>x"AF00",2858=>x"AF00",2859=>x"AF00",
2860=>x"AF00",2861=>x"AF00",2862=>x"AF00",2863=>x"AF00",2864=>x"AF00",
2865=>x"AF00",2866=>x"AF00",2867=>x"AF00",2868=>x"AF00",2869=>x"AF00",
2870=>x"AF00",2871=>x"AF00",2872=>x"AF00",2873=>x"AF00",2874=>x"AF00",
2875=>x"AF00",2876=>x"AF00",2877=>x"AF00",2878=>x"AF00",2879=>x"AF00",
2880=>x"AF00",2881=>x"AF00",2882=>x"AF00",2883=>x"AF00",2884=>x"AF00",
2885=>x"AF00",2886=>x"AF00",2887=>x"AF00",2888=>x"AF00",2889=>x"AF00",
2890=>x"AF00",2891=>x"AF00",2892=>x"AF00",2893=>x"AF00",2894=>x"AF00",
2895=>x"AF00",2896=>x"AF00",2897=>x"AF00",2898=>x"AF00",2899=>x"AF00",
2900=>x"AF00",2901=>x"AF00",2902=>x"AF00",2903=>x"AF00",2904=>x"AF00",
2905=>x"AF00",2906=>x"AF00",2907=>x"AF00",2908=>x"AF00",2909=>x"AF00",
2910=>x"AF00",2911=>x"AF00",2912=>x"AF00",2913=>x"AF00",2914=>x"AF00",
2915=>x"AF00",2916=>x"AF00",2917=>x"AF00",2918=>x"AF00",2919=>x"AF00",
2920=>x"AF00",2921=>x"AF00",2922=>x"AF00",2923=>x"AF00",2924=>x"AF00",
2925=>x"AF00",2926=>x"AF00",2927=>x"AF00",2928=>x"AF00",2929=>x"AF00",
2930=>x"AF00",2931=>x"AF00",2932=>x"AF00",2933=>x"AF00",2934=>x"AF00",
2935=>x"AF00",2936=>x"AF00",2937=>x"AF00",2938=>x"AF00",2939=>x"AF00",
2940=>x"AF00",2941=>x"AF00",2942=>x"AF00",2943=>x"AF00",2944=>x"AF00",
2945=>x"AF00",2946=>x"AF00",2947=>x"AF00",2948=>x"AF00",2949=>x"AF00",
2950=>x"AF00",2951=>x"AF00",2952=>x"AF00",2953=>x"AF00",2954=>x"AF00",
2955=>x"AF00",2956=>x"AF00",2957=>x"AF00",2958=>x"AF00",2959=>x"AF00",
2960=>x"AF00",2961=>x"AF00",2962=>x"AF00",2963=>x"AF00",2964=>x"AF00",
2965=>x"AF00",2966=>x"AF00",2967=>x"AF00",2968=>x"AF00",2969=>x"AF00",
2970=>x"AF00",2971=>x"AF00",2972=>x"AF00",2973=>x"AF00",2974=>x"AF00",
2975=>x"AF00",2976=>x"AF00",2977=>x"AF00",2978=>x"AF00",2979=>x"AF00",
2980=>x"AF00",2981=>x"AF00",2982=>x"AF00",2983=>x"AF00",2984=>x"AF00",
2985=>x"AF00",2986=>x"AF00",2987=>x"AF00",2988=>x"AF00",2989=>x"AF00",
2990=>x"AF00",2991=>x"AF00",2992=>x"AF00",2993=>x"AF00",2994=>x"AF00",
2995=>x"AF00",2996=>x"AF00",2997=>x"AF00",2998=>x"AF00",2999=>x"AF00",
3000=>x"AF00",3001=>x"AF00",3002=>x"AF00",3003=>x"AF00",3004=>x"AF00",
3005=>x"AF00",3006=>x"AF00",3007=>x"AF00",3008=>x"AF00",3009=>x"AF00",
3010=>x"AF00",3011=>x"AF00",3012=>x"AF00",3013=>x"AF00",3014=>x"AF00",
3015=>x"AF00",3016=>x"AF00",3017=>x"AF00",3018=>x"AF00",3019=>x"AF00",
3020=>x"AF00",3021=>x"AF00",3022=>x"AF00",3023=>x"AF00",3024=>x"AF00",
3025=>x"AF00",3026=>x"AF00",3027=>x"AF00",3028=>x"AF00",3029=>x"AF00",
3030=>x"AF00",3031=>x"AF00",3032=>x"AF00",3033=>x"AF00",3034=>x"AF00",
3035=>x"AF00",3036=>x"AF00",3037=>x"AF00",3038=>x"AF00",3039=>x"AF00",
3040=>x"AF00",3041=>x"AF00",3042=>x"AF00",3043=>x"AF00",3044=>x"AF00",
3045=>x"AF00",3046=>x"AF00",3047=>x"AF00",3048=>x"AF00",3049=>x"AF00",
3050=>x"AF00",3051=>x"AF00",3052=>x"AF00",3053=>x"AF00",3054=>x"AF00",
3055=>x"AF00",3056=>x"AF00",3057=>x"AF00",3058=>x"AF00",3059=>x"AF00",
3060=>x"AF00",3061=>x"AF00",3062=>x"AF00",3063=>x"AF00",3064=>x"AF00",
3065=>x"AF00",3066=>x"AF00",3067=>x"AF00",3068=>x"AF00",3069=>x"AF00",
3070=>x"AF00",3071=>x"AF00",3072=>x"AF00",3073=>x"AF00",3074=>x"AF00",
3075=>x"AF00",3076=>x"AF00",3077=>x"AF00",3078=>x"AF00",3079=>x"AF00",
3080=>x"AF00",3081=>x"AF00",3082=>x"AF00",3083=>x"AF00",3084=>x"AF00",
3085=>x"AF00",3086=>x"AF00",3087=>x"AF00",3088=>x"AF00",3089=>x"AF00",
3090=>x"AF00",3091=>x"AF00",3092=>x"AF00",3093=>x"AF00",3094=>x"AF00",
3095=>x"AF00",3096=>x"AF00",3097=>x"AF00",3098=>x"AF00",3099=>x"AF00",
3100=>x"AF00",3101=>x"AF00",3102=>x"AF00",3103=>x"AF00",3104=>x"AF00",
3105=>x"AF00",3106=>x"AF00",3107=>x"AF00",3108=>x"AF00",3109=>x"AF00",
3110=>x"AF00",3111=>x"AF00",3112=>x"AF00",3113=>x"AF00",3114=>x"AF00",
3115=>x"AF00",3116=>x"AF00",3117=>x"AF00",3118=>x"AF00",3119=>x"AF00",
3120=>x"AF00",3121=>x"AF00",3122=>x"AF00",3123=>x"AF00",3124=>x"AF00",
3125=>x"AF00",3126=>x"AF00",3127=>x"AF00",3128=>x"AF00",3129=>x"AF00",
3130=>x"AF00",3131=>x"AF00",3132=>x"AF00",3133=>x"AF00",3134=>x"AF00",
3135=>x"AF00",3136=>x"AF00",3137=>x"AF00",3138=>x"AF00",3139=>x"AF00",
3140=>x"AF00",3141=>x"AF00",3142=>x"AF00",3143=>x"AF00",3144=>x"AF00",
3145=>x"AF00",3146=>x"AF00",3147=>x"AF00",3148=>x"AF00",3149=>x"AF00",
3150=>x"AF00",3151=>x"AF00",3152=>x"AF00",3153=>x"AF00",3154=>x"AF00",
3155=>x"AF00",3156=>x"AF00",3157=>x"AF00",3158=>x"AF00",3159=>x"AF00",
3160=>x"AF00",3161=>x"AF00",3162=>x"AF00",3163=>x"AF00",3164=>x"AF00",
3165=>x"AF00",3166=>x"AF00",3167=>x"AF00",3168=>x"AF00",3169=>x"AF00",
3170=>x"AF00",3171=>x"AF00",3172=>x"AF00",3173=>x"AF00",3174=>x"AF00",
3175=>x"AF00",3176=>x"AF00",3177=>x"AF00",3178=>x"AF00",3179=>x"AF00",
3180=>x"AF00",3181=>x"AF00",3182=>x"AF00",3183=>x"AF00",3184=>x"AF00",
3185=>x"AF00",3186=>x"AF00",3187=>x"AF00",3188=>x"AF00",3189=>x"AF00",
3190=>x"AF00",3191=>x"AF00",3192=>x"AF00",3193=>x"AF00",3194=>x"AF00",
3195=>x"AF00",3196=>x"AF00",3197=>x"AF00",3198=>x"AF00",3199=>x"AF00",
3200=>x"AF00",3201=>x"AF00",3202=>x"AF00",3203=>x"AF00",3204=>x"AF00",
3205=>x"AF00",3206=>x"AF00",3207=>x"AF00",3208=>x"AF00",3209=>x"AF00",
3210=>x"AF00",3211=>x"AF00",3212=>x"AF00",3213=>x"AF00",3214=>x"AF00",
3215=>x"AF00",3216=>x"AF00",3217=>x"AF00",3218=>x"AF00",3219=>x"AF00",
3220=>x"AF00",3221=>x"AF00",3222=>x"AF00",3223=>x"AF00",3224=>x"AF00",
3225=>x"AF00",3226=>x"AF00",3227=>x"AF00",3228=>x"AF00",3229=>x"AF00",
3230=>x"AF00",3231=>x"AF00",3232=>x"AF00",3233=>x"AF00",3234=>x"AF00",
3235=>x"AF00",3236=>x"AF00",3237=>x"AF00",3238=>x"AF00",3239=>x"AF00",
3240=>x"AF00",3241=>x"AF00",3242=>x"AF00",3243=>x"AF00",3244=>x"AF00",
3245=>x"AF00",3246=>x"AF00",3247=>x"AF00",3248=>x"AF00",3249=>x"AF00",
3250=>x"AF00",3251=>x"AF00",3252=>x"AF00",3253=>x"AF00",3254=>x"AF00",
3255=>x"AF00",3256=>x"AF00",3257=>x"AF00",3258=>x"AF00",3259=>x"AF00",
3260=>x"AF00",3261=>x"AF00",3262=>x"AF00",3263=>x"AF00",3264=>x"AF00",
3265=>x"AF00",3266=>x"AF00",3267=>x"AF00",3268=>x"AF00",3269=>x"AF00",
3270=>x"AF00",3271=>x"AF00",3272=>x"AF00",3273=>x"AF00",3274=>x"AF00",
3275=>x"AF00",3276=>x"AF00",3277=>x"AF00",3278=>x"AF00",3279=>x"AF00",
3280=>x"AF00",3281=>x"AF00",3282=>x"AF00",3283=>x"AF00",3284=>x"AF00",
3285=>x"AF00",3286=>x"AF00",3287=>x"AF00",3288=>x"AF00",3289=>x"AF00",
3290=>x"AF00",3291=>x"AF00",3292=>x"AF00",3293=>x"AF00",3294=>x"AF00",
3295=>x"AF00",3296=>x"AF00",3297=>x"AF00",3298=>x"AF00",3299=>x"AF00",
3300=>x"AF00",3301=>x"AF00",3302=>x"AF00",3303=>x"AF00",3304=>x"AF00",
3305=>x"AF00",3306=>x"AF00",3307=>x"AF00",3308=>x"AF00",3309=>x"AF00",
3310=>x"AF00",3311=>x"AF00",3312=>x"AF00",3313=>x"AF00",3314=>x"AF00",
3315=>x"AF00",3316=>x"AF00",3317=>x"AF00",3318=>x"AF00",3319=>x"AF00",
3320=>x"AF00",3321=>x"AF00",3322=>x"AF00",3323=>x"AF00",3324=>x"AF00",
3325=>x"AF00",3326=>x"AF00",3327=>x"AF00",3328=>x"AF00",3329=>x"AF00",
3330=>x"AF00",3331=>x"AF00",3332=>x"AF00",3333=>x"AF00",3334=>x"AF00",
3335=>x"AF00",3336=>x"AF00",3337=>x"AF00",3338=>x"AF00",3339=>x"AF00",
3340=>x"AF00",3341=>x"AF00",3342=>x"AF00",3343=>x"AF00",3344=>x"AF00",
3345=>x"AF00",3346=>x"AF00",3347=>x"AF00",3348=>x"AF00",3349=>x"AF00",
3350=>x"AF00",3351=>x"AF00",3352=>x"AF00",3353=>x"AF00",3354=>x"AF00",
3355=>x"AF00",3356=>x"AF00",3357=>x"AF00",3358=>x"AF00",3359=>x"AF00",
3360=>x"AF00",3361=>x"AF00",3362=>x"AF00",3363=>x"AF00",3364=>x"AF00",
3365=>x"AF00",3366=>x"AF00",3367=>x"AF00",3368=>x"AF00",3369=>x"AF00",
3370=>x"AF00",3371=>x"AF00",3372=>x"AF00",3373=>x"AF00",3374=>x"AF00",
3375=>x"AF00",3376=>x"AF00",3377=>x"AF00",3378=>x"AF00",3379=>x"AF00",
3380=>x"AF00",3381=>x"AF00",3382=>x"AF00",3383=>x"AF00",3384=>x"AF00",
3385=>x"AF00",3386=>x"AF00",3387=>x"AF00",3388=>x"AF00",3389=>x"AF00",
3390=>x"AF00",3391=>x"AF00",3392=>x"AF00",3393=>x"AF00",3394=>x"AF00",
3395=>x"AF00",3396=>x"AF00",3397=>x"AF00",3398=>x"AF00",3399=>x"AF00",
3400=>x"AF00",3401=>x"AF00",3402=>x"AF00",3403=>x"AF00",3404=>x"AF00",
3405=>x"AF00",3406=>x"AF00",3407=>x"AF00",3408=>x"AF00",3409=>x"AF00",
3410=>x"AF00",3411=>x"AF00",3412=>x"AF00",3413=>x"AF00",3414=>x"AF00",
3415=>x"AF00",3416=>x"AF00",3417=>x"AF00",3418=>x"AF00",3419=>x"AF00",
3420=>x"AF00",3421=>x"AF00",3422=>x"AF00",3423=>x"AF00",3424=>x"AF00",
3425=>x"AF00",3426=>x"AF00",3427=>x"AF00",3428=>x"AF00",3429=>x"AF00",
3430=>x"AF00",3431=>x"AF00",3432=>x"AF00",3433=>x"AF00",3434=>x"AF00",
3435=>x"AF00",3436=>x"AF00",3437=>x"AF00",3438=>x"AF00",3439=>x"AF00",
3440=>x"AF00",3441=>x"AF00",3442=>x"AF00",3443=>x"AF00",3444=>x"AF00",
3445=>x"AF00",3446=>x"AF00",3447=>x"AF00",3448=>x"AF00",3449=>x"AF00",
3450=>x"AF00",3451=>x"AF00",3452=>x"AF00",3453=>x"AF00",3454=>x"AF00",
3455=>x"AF00",3456=>x"AF00",3457=>x"AF00",3458=>x"AF00",3459=>x"AF00",
3460=>x"AF00",3461=>x"AF00",3462=>x"AF00",3463=>x"AF00",3464=>x"AF00",
3465=>x"AF00",3466=>x"AF00",3467=>x"AF00",3468=>x"AF00",3469=>x"AF00",
3470=>x"AF00",3471=>x"AF00",3472=>x"AF00",3473=>x"AF00",3474=>x"AF00",
3475=>x"AF00",3476=>x"AF00",3477=>x"AF00",3478=>x"AF00",3479=>x"AF00",
3480=>x"AF00",3481=>x"AF00",3482=>x"AF00",3483=>x"AF00",3484=>x"AF00",
3485=>x"AF00",3486=>x"AF00",3487=>x"AF00",3488=>x"AF00",3489=>x"AF00",
3490=>x"AF00",3491=>x"AF00",3492=>x"AF00",3493=>x"AF00",3494=>x"AF00",
3495=>x"AF00",3496=>x"AF00",3497=>x"AF00",3498=>x"AF00",3499=>x"AF00",
3500=>x"AF00",3501=>x"AF00",3502=>x"AF00",3503=>x"AF00",3504=>x"AF00",
3505=>x"AF00",3506=>x"AF00",3507=>x"AF00",3508=>x"AF00",3509=>x"AF00",
3510=>x"AF00",3511=>x"AF00",3512=>x"AF00",3513=>x"AF00",3514=>x"AF00",
3515=>x"AF00",3516=>x"AF00",3517=>x"AF00",3518=>x"AF00",3519=>x"AF00",
3520=>x"AF00",3521=>x"AF00",3522=>x"AF00",3523=>x"AF00",3524=>x"AF00",
3525=>x"AF00",3526=>x"AF00",3527=>x"AF00",3528=>x"AF00",3529=>x"AF00",
3530=>x"AF00",3531=>x"AF00",3532=>x"AF00",3533=>x"AF00",3534=>x"AF00",
3535=>x"AF00",3536=>x"AF00",3537=>x"AF00",3538=>x"AF00",3539=>x"AF00",
3540=>x"AF00",3541=>x"AF00",3542=>x"AF00",3543=>x"AF00",3544=>x"AF00",
3545=>x"AF00",3546=>x"AF00",3547=>x"AF00",3548=>x"AF00",3549=>x"AF00",
3550=>x"AF00",3551=>x"AF00",3552=>x"AF00",3553=>x"AF00",3554=>x"AF00",
3555=>x"AF00",3556=>x"AF00",3557=>x"AF00",3558=>x"AF00",3559=>x"AF00",
3560=>x"AF00",3561=>x"AF00",3562=>x"AF00",3563=>x"AF00",3564=>x"AF00",
3565=>x"AF00",3566=>x"AF00",3567=>x"AF00",3568=>x"AF00",3569=>x"AF00",
3570=>x"AF00",3571=>x"AF00",3572=>x"AF00",3573=>x"AF00",3574=>x"AF00",
3575=>x"AF00",3576=>x"AF00",3577=>x"AF00",3578=>x"AF00",3579=>x"AF00",
3580=>x"AF00",3581=>x"AF00",3582=>x"AF00",3583=>x"AF00",3584=>x"AF00",
3585=>x"AF00",3586=>x"AF00",3587=>x"AF00",3588=>x"AF00",3589=>x"AF00",
3590=>x"AF00",3591=>x"AF00",3592=>x"AF00",3593=>x"AF00",3594=>x"AF00",
3595=>x"AF00",3596=>x"AF00",3597=>x"AF00",3598=>x"AF00",3599=>x"AF00",
3600=>x"AF00",3601=>x"AF00",3602=>x"AF00",3603=>x"AF00",3604=>x"AF00",
3605=>x"AF00",3606=>x"AF00",3607=>x"AF00",3608=>x"AF00",3609=>x"AF00",
3610=>x"AF00",3611=>x"AF00",3612=>x"AF00",3613=>x"AF00",3614=>x"AF00",
3615=>x"AF00",3616=>x"AF00",3617=>x"AF00",3618=>x"AF00",3619=>x"AF00",
3620=>x"AF00",3621=>x"AF00",3622=>x"AF00",3623=>x"AF00",3624=>x"AF00",
3625=>x"AF00",3626=>x"AF00",3627=>x"AF00",3628=>x"AF00",3629=>x"AF00",
3630=>x"AF00",3631=>x"AF00",3632=>x"AF00",3633=>x"AF00",3634=>x"AF00",
3635=>x"AF00",3636=>x"AF00",3637=>x"AF00",3638=>x"AF00",3639=>x"AF00",
3640=>x"AF00",3641=>x"AF00",3642=>x"AF00",3643=>x"AF00",3644=>x"AF00",
3645=>x"AF00",3646=>x"AF00",3647=>x"AF00",3648=>x"AF00",3649=>x"AF00",
3650=>x"AF00",3651=>x"AF00",3652=>x"AF00",3653=>x"AF00",3654=>x"AF00",
3655=>x"AF00",3656=>x"AF00",3657=>x"AF00",3658=>x"AF00",3659=>x"AF00",
3660=>x"AF00",3661=>x"AF00",3662=>x"AF00",3663=>x"AF00",3664=>x"AF00",
3665=>x"AF00",3666=>x"AF00",3667=>x"AF00",3668=>x"AF00",3669=>x"AF00",
3670=>x"AF00",3671=>x"AF00",3672=>x"AF00",3673=>x"AF00",3674=>x"AF00",
3675=>x"AF00",3676=>x"AF00",3677=>x"AF00",3678=>x"AF00",3679=>x"AF00",
3680=>x"AF00",3681=>x"AF00",3682=>x"AF00",3683=>x"AF00",3684=>x"AF00",
3685=>x"AF00",3686=>x"AF00",3687=>x"AF00",3688=>x"AF00",3689=>x"AF00",
3690=>x"AF00",3691=>x"AF00",3692=>x"AF00",3693=>x"AF00",3694=>x"AF00",
3695=>x"AF00",3696=>x"AF00",3697=>x"AF00",3698=>x"AF00",3699=>x"AF00",
3700=>x"AF00",3701=>x"AF00",3702=>x"AF00",3703=>x"AF00",3704=>x"AF00",
3705=>x"AF00",3706=>x"AF00",3707=>x"AF00",3708=>x"AF00",3709=>x"AF00",
3710=>x"AF00",3711=>x"AF00",3712=>x"AF00",3713=>x"AF00",3714=>x"AF00",
3715=>x"AF00",3716=>x"AF00",3717=>x"AF00",3718=>x"AF00",3719=>x"AF00",
3720=>x"AF00",3721=>x"AF00",3722=>x"AF00",3723=>x"AF00",3724=>x"AF00",
3725=>x"AF00",3726=>x"AF00",3727=>x"AF00",3728=>x"AF00",3729=>x"AF00",
3730=>x"AF00",3731=>x"AF00",3732=>x"AF00",3733=>x"AF00",3734=>x"AF00",
3735=>x"AF00",3736=>x"AF00",3737=>x"AF00",3738=>x"AF00",3739=>x"AF00",
3740=>x"AF00",3741=>x"AF00",3742=>x"AF00",3743=>x"AF00",3744=>x"AF00",
3745=>x"AF00",3746=>x"AF00",3747=>x"AF00",3748=>x"AF00",3749=>x"AF00",
3750=>x"AF00",3751=>x"AF00",3752=>x"AF00",3753=>x"AF00",3754=>x"AF00",
3755=>x"AF00",3756=>x"AF00",3757=>x"AF00",3758=>x"AF00",3759=>x"AF00",
3760=>x"AF00",3761=>x"AF00",3762=>x"AF00",3763=>x"AF00",3764=>x"AF00",
3765=>x"AF00",3766=>x"AF00",3767=>x"AF00",3768=>x"AF00",3769=>x"AF00",
3770=>x"AF00",3771=>x"AF00",3772=>x"AF00",3773=>x"AF00",3774=>x"AF00",
3775=>x"AF00",3776=>x"AF00",3777=>x"AF00",3778=>x"AF00",3779=>x"AF00",
3780=>x"AF00",3781=>x"AF00",3782=>x"AF00",3783=>x"AF00",3784=>x"AF00",
3785=>x"AF00",3786=>x"AF00",3787=>x"AF00",3788=>x"AF00",3789=>x"AF00",
3790=>x"AF00",3791=>x"AF00",3792=>x"AF00",3793=>x"AF00",3794=>x"AF00",
3795=>x"AF00",3796=>x"AF00",3797=>x"AF00",3798=>x"AF00",3799=>x"AF00",
3800=>x"AF00",3801=>x"AF00",3802=>x"AF00",3803=>x"AF00",3804=>x"AF00",
3805=>x"AF00",3806=>x"AF00",3807=>x"AF00",3808=>x"AF00",3809=>x"AF00",
3810=>x"AF00",3811=>x"AF00",3812=>x"AF00",3813=>x"AF00",3814=>x"AF00",
3815=>x"AF00",3816=>x"AF00",3817=>x"AF00",3818=>x"AF00",3819=>x"AF00",
3820=>x"AF00",3821=>x"AF00",3822=>x"AF00",3823=>x"AF00",3824=>x"AF00",
3825=>x"AF00",3826=>x"AF00",3827=>x"AF00",3828=>x"AF00",3829=>x"AF00",
3830=>x"AF00",3831=>x"AF00",3832=>x"AF00",3833=>x"AF00",3834=>x"AF00",
3835=>x"AF00",3836=>x"AF00",3837=>x"AF00",3838=>x"AF00",3839=>x"AF00",
3840=>x"AF00",3841=>x"AF00",3842=>x"AF00",3843=>x"AF00",3844=>x"AF00",
3845=>x"AF00",3846=>x"AF00",3847=>x"AF00",3848=>x"AF00",3849=>x"AF00",
3850=>x"AF00",3851=>x"AF00",3852=>x"AF00",3853=>x"AF00",3854=>x"AF00",
3855=>x"AF00",3856=>x"AF00",3857=>x"AF00",3858=>x"AF00",3859=>x"AF00",
3860=>x"AF00",3861=>x"AF00",3862=>x"AF00",3863=>x"AF00",3864=>x"AF00",
3865=>x"AF00",3866=>x"AF00",3867=>x"AF00",3868=>x"AF00",3869=>x"AF00",
3870=>x"AF00",3871=>x"AF00",3872=>x"AF00",3873=>x"AF00",3874=>x"AF00",
3875=>x"AF00",3876=>x"AF00",3877=>x"AF00",3878=>x"AF00",3879=>x"AF00",
3880=>x"AF00",3881=>x"AF00",3882=>x"AF00",3883=>x"AF00",3884=>x"AF00",
3885=>x"AF00",3886=>x"AF00",3887=>x"AF00",3888=>x"AF00",3889=>x"AF00",
3890=>x"AF00",3891=>x"AF00",3892=>x"AF00",3893=>x"AF00",3894=>x"AF00",
3895=>x"AF00",3896=>x"AF00",3897=>x"AF00",3898=>x"AF00",3899=>x"AF00",
3900=>x"AF00",3901=>x"AF00",3902=>x"AF00",3903=>x"AF00",3904=>x"AF00",
3905=>x"AF00",3906=>x"AF00",3907=>x"AF00",3908=>x"AF00",3909=>x"AF00",
3910=>x"AF00",3911=>x"AF00",3912=>x"AF00",3913=>x"AF00",3914=>x"AF00",
3915=>x"AF00",3916=>x"AF00",3917=>x"AF00",3918=>x"AF00",3919=>x"AF00",
3920=>x"AF00",3921=>x"AF00",3922=>x"AF00",3923=>x"AF00",3924=>x"AF00",
3925=>x"AF00",3926=>x"AF00",3927=>x"AF00",3928=>x"AF00",3929=>x"AF00",
3930=>x"AF00",3931=>x"AF00",3932=>x"AF00",3933=>x"AF00",3934=>x"AF00",
3935=>x"AF00",3936=>x"AF00",3937=>x"AF00",3938=>x"AF00",3939=>x"AF00",
3940=>x"AF00",3941=>x"AF00",3942=>x"AF00",3943=>x"AF00",3944=>x"AF00",
3945=>x"AF00",3946=>x"AF00",3947=>x"AF00",3948=>x"AF00",3949=>x"AF00",
3950=>x"AF00",3951=>x"AF00",3952=>x"AF00",3953=>x"AF00",3954=>x"AF00",
3955=>x"AF00",3956=>x"AF00",3957=>x"AF00",3958=>x"AF00",3959=>x"AF00",
3960=>x"AF00",3961=>x"AF00",3962=>x"AF00",3963=>x"AF00",3964=>x"AF00",
3965=>x"AF00",3966=>x"AF00",3967=>x"AF00",3968=>x"AF00",3969=>x"AF00",
3970=>x"AF00",3971=>x"AF00",3972=>x"AF00",3973=>x"AF00",3974=>x"AF00",
3975=>x"AF00",3976=>x"AF00",3977=>x"AF00",3978=>x"AF00",3979=>x"AF00",
3980=>x"AF00",3981=>x"AF00",3982=>x"AF00",3983=>x"AF00",3984=>x"AF00",
3985=>x"AF00",3986=>x"AF00",3987=>x"AF00",3988=>x"AF00",3989=>x"AF00",
3990=>x"AF00",3991=>x"AF00",3992=>x"AF00",3993=>x"AF00",3994=>x"AF00",
3995=>x"AF00",3996=>x"AF00",3997=>x"AF00",3998=>x"AF00",3999=>x"AF00",
4000=>x"AF00",4001=>x"AF00",4002=>x"AF00",4003=>x"AF00",4004=>x"AF00",
4005=>x"AF00",4006=>x"AF00",4007=>x"AF00",4008=>x"AF00",4009=>x"AF00",
4010=>x"AF00",4011=>x"AF00",4012=>x"AF00",4013=>x"AF00",4014=>x"AF00",
4015=>x"AF00",4016=>x"AF00",4017=>x"AF00",4018=>x"AF00",4019=>x"AF00",
4020=>x"AF00",4021=>x"AF00",4022=>x"AF00",4023=>x"AF00",4024=>x"AF00",
4025=>x"AF00",4026=>x"AF00",4027=>x"AF00",4028=>x"AF00",4029=>x"AF00",
4030=>x"AF00",4031=>x"AF00",4032=>x"AF00",4033=>x"AF00",4034=>x"AF00",
4035=>x"AF00",4036=>x"AF00",4037=>x"AF00",4038=>x"AF00",4039=>x"AF00",
4040=>x"AF00",4041=>x"AF00",4042=>x"AF00",4043=>x"AF00",4044=>x"AF00",
4045=>x"AF00",4046=>x"AF00",4047=>x"AF00",4048=>x"AF00",4049=>x"AF00",
4050=>x"AF00",4051=>x"AF00",4052=>x"AF00",4053=>x"AF00",4054=>x"AF00",
4055=>x"AF00",4056=>x"AF00",4057=>x"AF00",4058=>x"AF00",4059=>x"AF00",
4060=>x"AF00",4061=>x"AF00",4062=>x"AF00",4063=>x"AF00",4064=>x"AF00",
4065=>x"AF00",4066=>x"AF00",4067=>x"AF00",4068=>x"AF00",4069=>x"AF00",
4070=>x"AF00",4071=>x"AF00",4072=>x"AF00",4073=>x"AF00",4074=>x"AF00",
4075=>x"AF00",4076=>x"AF00",4077=>x"AF00",4078=>x"AF00",4079=>x"AF00",
4080=>x"AF00",4081=>x"AF00",4082=>x"AF00",4083=>x"AF00",4084=>x"AF00",
4085=>x"AF00",4086=>x"AF00",4087=>x"AF00",4088=>x"AF00",4089=>x"AF00",
4090=>x"AF00",4091=>x"AF00",4092=>x"A008",4093=>x"0F1F",4094=>x"A02E",
4095=>x"A002",4096=>x"0110",4097=>x"C822",4098=>x"2FD3",4099=>x"A0F8",
4100=>x"48E0",4101=>x"0801",4102=>x"AF00",4103=>x"AF00",4104=>x"AF00",
4105=>x"AF00",4106=>x"AF00",4107=>x"AF00",4108=>x"AF00",4109=>x"AF00",
4110=>x"AF00",4111=>x"AF00",4112=>x"AF00",4113=>x"AF00",4114=>x"AF00",
4115=>x"AF00",4116=>x"AF00",4117=>x"AF00",4118=>x"AF00",4119=>x"AF00",
4120=>x"AF00",4121=>x"AF00",4122=>x"AF00",4123=>x"AF00",4124=>x"AF00",
4125=>x"AF00",4126=>x"AF00",4127=>x"AF00",4128=>x"AF00",4129=>x"AF00",
4130=>x"AF00",4131=>x"AF00",4132=>x"AF00",4133=>x"AF00",4134=>x"AF00",
4135=>x"AF00",4136=>x"AF00",4137=>x"AF00",4138=>x"AF00",4139=>x"AF00",
4140=>x"AF00",4141=>x"AF00",4142=>x"AF00",4143=>x"AF00",4144=>x"AF00",
4145=>x"AF00",4146=>x"AF00",4147=>x"AF00",4148=>x"AF00",4149=>x"AF00",
4150=>x"AF00",4151=>x"AF00",4152=>x"AF00",4153=>x"AF00",4154=>x"AF00",
4155=>x"AF00",4156=>x"AF00",4157=>x"AF00",4158=>x"AF00",4159=>x"AF00",
4160=>x"AF00",4161=>x"AF00",4162=>x"AF00",4163=>x"AF00",4164=>x"AF00",
4165=>x"AF00",4166=>x"AF00",4167=>x"AF00",4168=>x"AF00",4169=>x"AF00",
4170=>x"AF00",4171=>x"AF00",4172=>x"AF00",4173=>x"AF00",4174=>x"AF00",
4175=>x"AF00",4176=>x"AF00",4177=>x"AF00",4178=>x"AF00",4179=>x"AF00",
4180=>x"AF00",4181=>x"AF00",4182=>x"AF00",4183=>x"AF00",4184=>x"AF00",
4185=>x"AF00",4186=>x"AF00",4187=>x"AF00",4188=>x"AF00",4189=>x"AF00",
4190=>x"AF00",4191=>x"AF00",4192=>x"AF00",4193=>x"AF00",4194=>x"AF00",
4195=>x"AF00",4196=>x"AF00",4197=>x"AF00",4198=>x"AF00",4199=>x"AF00",
4200=>x"AF00",4201=>x"AF00",4202=>x"AF00",4203=>x"AF00",4204=>x"AF00",
4205=>x"AF00",4206=>x"AF00",4207=>x"AF00",4208=>x"AF00",4209=>x"AF00",
4210=>x"AF00",4211=>x"AF00",4212=>x"AF00",4213=>x"AF00",4214=>x"AF00",
4215=>x"AF00",4216=>x"AF00",4217=>x"AF00",4218=>x"AF00",4219=>x"AF00",
4220=>x"AF00",4221=>x"AF00",4222=>x"AF00",4223=>x"AF00",4224=>x"AF00",
4225=>x"AF00",4226=>x"AF00",4227=>x"AF00",4228=>x"AF00",4229=>x"AF00",
4230=>x"AF00",4231=>x"AF00",4232=>x"AF00",4233=>x"AF00",4234=>x"AF00",
4235=>x"AF00",4236=>x"AF00",4237=>x"AF00",4238=>x"AF00",4239=>x"AF00",
4240=>x"AF00",4241=>x"AF00",4242=>x"AF00",4243=>x"AF00",4244=>x"AF00",
4245=>x"AF00",4246=>x"AF00",4247=>x"AF00",4248=>x"AF00",4249=>x"AF00",
4250=>x"AF00",4251=>x"AF00",4252=>x"AF00",4253=>x"AF00",4254=>x"AF00",
4255=>x"AF00",4256=>x"AF00",4257=>x"AF00",4258=>x"AF00",4259=>x"AF00",
4260=>x"AF00",4261=>x"AF00",4262=>x"AF00",4263=>x"AF00",4264=>x"AF00",
4265=>x"AF00",4266=>x"AF00",4267=>x"AF00",4268=>x"AF00",4269=>x"AF00",
4270=>x"AF00",4271=>x"AF00",4272=>x"AF00",4273=>x"AF00",4274=>x"AF00",
4275=>x"AF00",4276=>x"AF00",4277=>x"AF00",4278=>x"AF00",4279=>x"AF00",
4280=>x"AF00",4281=>x"AF00",4282=>x"AF00",4283=>x"AF00",4284=>x"AF00",
4285=>x"AF00",4286=>x"AF00",4287=>x"AF00",4288=>x"AF00",4289=>x"AF00",
4290=>x"AF00",4291=>x"AF00",4292=>x"AF00",4293=>x"AF00",4294=>x"AF00",
4295=>x"AF00",4296=>x"AF00",4297=>x"AF00",4298=>x"AF00",4299=>x"AF00",
4300=>x"AF00",4301=>x"AF00",4302=>x"AF00",4303=>x"AF00",4304=>x"AF00",
4305=>x"AF00",4306=>x"AF00",4307=>x"AF00",4308=>x"AF00",4309=>x"AF00",
4310=>x"AF00",4311=>x"AF00",4312=>x"AF00",4313=>x"AF00",4314=>x"AF00",
4315=>x"AF00",4316=>x"AF00",4317=>x"AF00",4318=>x"AF00",4319=>x"AF00",
4320=>x"AF00",4321=>x"AF00",4322=>x"AF00",4323=>x"AF00",4324=>x"AF00",
4325=>x"AF00",4326=>x"AF00",4327=>x"AF00",4328=>x"AF00",4329=>x"AF00",
4330=>x"AF00",4331=>x"AF00",4332=>x"AF00",4333=>x"AF00",4334=>x"AF00",
4335=>x"AF00",4336=>x"AF00",4337=>x"AF00",4338=>x"AF00",4339=>x"AF00",
4340=>x"AF00",4341=>x"AF00",4342=>x"AF00",4343=>x"AF00",4344=>x"AF00",
4345=>x"AF00",4346=>x"AF00",4347=>x"AF00",4348=>x"AF00",4349=>x"AF00",
4350=>x"AF00",4351=>x"AF00",4352=>x"AF00",4353=>x"AF00",4354=>x"AF00",
4355=>x"AF00",4356=>x"AF00",4357=>x"AF00",4358=>x"AF00",4359=>x"AF00",
4360=>x"AF00",4361=>x"AF00",4362=>x"AF00",4363=>x"AF00",4364=>x"AF00",
4365=>x"AF00",4366=>x"AF00",4367=>x"AF00",4368=>x"AF00",4369=>x"AF00",
4370=>x"AF00",4371=>x"AF00",4372=>x"AF00",4373=>x"AF00",4374=>x"AF00",
4375=>x"AF00",4376=>x"AF00",4377=>x"AF00",4378=>x"AF00",4379=>x"AF00",
4380=>x"AF00",4381=>x"AF00",4382=>x"AF00",4383=>x"AF00",4384=>x"AF00",
4385=>x"AF00",4386=>x"AF00",4387=>x"AF00",4388=>x"AF00",4389=>x"AF00",
4390=>x"AF00",4391=>x"AF00",4392=>x"AF00",4393=>x"AF00",4394=>x"AF00",
4395=>x"AF00",4396=>x"AF00",4397=>x"AF00",4398=>x"AF00",4399=>x"AF00",
4400=>x"AF00",4401=>x"AF00",4402=>x"AF00",4403=>x"AF00",4404=>x"AF00",
4405=>x"AF00",4406=>x"AF00",4407=>x"AF00",4408=>x"AF00",4409=>x"AF00",
4410=>x"AF00",4411=>x"AF00",4412=>x"AF00",4413=>x"AF00",4414=>x"AF00",
4415=>x"AF00",4416=>x"AF00",4417=>x"AF00",4418=>x"AF00",4419=>x"AF00",
4420=>x"AF00",4421=>x"AF00",4422=>x"AF00",4423=>x"AF00",4424=>x"AF00",
4425=>x"AF00",4426=>x"AF00",4427=>x"AF00",4428=>x"AF00",4429=>x"AF00",
4430=>x"AF00",4431=>x"AF00",4432=>x"AF00",4433=>x"AF00",4434=>x"AF00",
4435=>x"AF00",4436=>x"AF00",4437=>x"AF00",4438=>x"AF00",4439=>x"AF00",
4440=>x"AF00",4441=>x"AF00",4442=>x"AF00",4443=>x"AF00",4444=>x"AF00",
4445=>x"AF00",4446=>x"AF00",4447=>x"AF00",4448=>x"AF00",4449=>x"AF00",
4450=>x"AF00",4451=>x"AF00",4452=>x"AF00",4453=>x"AF00",4454=>x"AF00",
4455=>x"AF00",4456=>x"AF00",4457=>x"AF00",4458=>x"AF00",4459=>x"AF00",
4460=>x"AF00",4461=>x"AF00",4462=>x"AF00",4463=>x"AF00",4464=>x"AF00",
4465=>x"AF00",4466=>x"AF00",4467=>x"AF00",4468=>x"AF00",4469=>x"AF00",
4470=>x"AF00",4471=>x"AF00",4472=>x"AF00",4473=>x"AF00",4474=>x"AF00",
4475=>x"AF00",4476=>x"AF00",4477=>x"AF00",4478=>x"AF00",4479=>x"AF00",
4480=>x"AF00",4481=>x"AF00",4482=>x"AF00",4483=>x"AF00",4484=>x"AF00",
4485=>x"AF00",4486=>x"AF00",4487=>x"AF00",4488=>x"AF00",4489=>x"AF00",
4490=>x"AF00",4491=>x"AF00",4492=>x"AF00",4493=>x"AF00",4494=>x"AF00",
4495=>x"AF00",4496=>x"AF00",4497=>x"AF00",4498=>x"AF00",4499=>x"AF00",
4500=>x"AF00",4501=>x"AF00",4502=>x"AF00",4503=>x"AF00",4504=>x"AF00",
4505=>x"AF00",4506=>x"AF00",4507=>x"AF00",4508=>x"AF00",4509=>x"AF00",
4510=>x"AF00",4511=>x"AF00",4512=>x"AF00",4513=>x"AF00",4514=>x"AF00",
4515=>x"AF00",4516=>x"AF00",4517=>x"AF00",4518=>x"AF00",4519=>x"AF00",
4520=>x"AF00",4521=>x"AF00",4522=>x"AF00",4523=>x"AF00",4524=>x"AF00",
4525=>x"AF00",4526=>x"AF00",4527=>x"AF00",4528=>x"AF00",4529=>x"AF00",
4530=>x"AF00",4531=>x"AF00",4532=>x"AF00",4533=>x"AF00",4534=>x"AF00",
4535=>x"AF00",4536=>x"AF00",4537=>x"AF00",4538=>x"AF00",4539=>x"AF00",
4540=>x"AF00",4541=>x"AF00",4542=>x"AF00",4543=>x"AF00",4544=>x"AF00",
4545=>x"AF00",4546=>x"AF00",4547=>x"AF00",4548=>x"AF00",4549=>x"AF00",
4550=>x"AF00",4551=>x"AF00",4552=>x"AF00",4553=>x"AF00",4554=>x"AF00",
4555=>x"AF00",4556=>x"AF00",4557=>x"AF00",4558=>x"AF00",4559=>x"AF00",
4560=>x"AF00",4561=>x"AF00",4562=>x"AF00",4563=>x"AF00",4564=>x"AF00",
4565=>x"AF00",4566=>x"AF00",4567=>x"AF00",4568=>x"AF00",4569=>x"AF00",
4570=>x"AF00",4571=>x"AF00",4572=>x"AF00",4573=>x"AF00",4574=>x"AF00",
4575=>x"AF00",4576=>x"AF00",4577=>x"AF00",4578=>x"AF00",4579=>x"AF00",
4580=>x"AF00",4581=>x"AF00",4582=>x"AF00",4583=>x"AF00",4584=>x"AF00",
4585=>x"AF00",4586=>x"AF00",4587=>x"AF00",4588=>x"AF00",4589=>x"AF00",
4590=>x"AF00",4591=>x"AF00",4592=>x"AF00",4593=>x"AF00",4594=>x"AF00",
4595=>x"AF00",4596=>x"AF00",4597=>x"AF00",4598=>x"AF00",4599=>x"AF00",
4600=>x"AF00",4601=>x"AF00",4602=>x"AF00",4603=>x"AF00",4604=>x"AF00",
4605=>x"AF00",4606=>x"AF00",4607=>x"AF00",4608=>x"AF00",4609=>x"AF00",
4610=>x"AF00",4611=>x"AF00",4612=>x"AF00",4613=>x"AF00",4614=>x"AF00",
4615=>x"AF00",4616=>x"AF00",4617=>x"AF00",4618=>x"AF00",4619=>x"AF00",
4620=>x"AF00",4621=>x"AF00",4622=>x"AF00",4623=>x"AF00",4624=>x"AF00",
4625=>x"AF00",4626=>x"AF00",4627=>x"AF00",4628=>x"AF00",4629=>x"AF00",
4630=>x"AF00",4631=>x"AF00",4632=>x"AF00",4633=>x"AF00",4634=>x"AF00",
4635=>x"AF00",4636=>x"AF00",4637=>x"AF00",4638=>x"AF00",4639=>x"AF00",
4640=>x"AF00",4641=>x"AF00",4642=>x"AF00",4643=>x"AF00",4644=>x"AF00",
4645=>x"AF00",4646=>x"AF00",4647=>x"AF00",4648=>x"AF00",4649=>x"AF00",
4650=>x"AF00",4651=>x"AF00",4652=>x"AF00",4653=>x"AF00",4654=>x"AF00",
4655=>x"AF00",4656=>x"AF00",4657=>x"AF00",4658=>x"AF00",4659=>x"AF00",
4660=>x"AF00",4661=>x"AF00",4662=>x"AF00",4663=>x"AF00",4664=>x"AF00",
4665=>x"AF00",4666=>x"AF00",4667=>x"AF00",4668=>x"AF00",4669=>x"AF00",
4670=>x"AF00",4671=>x"AF00",4672=>x"AF00",4673=>x"AF00",4674=>x"AF00",
4675=>x"AF00",4676=>x"AF00",4677=>x"AF00",4678=>x"AF00",4679=>x"AF00",
4680=>x"AF00",4681=>x"AF00",4682=>x"AF00",4683=>x"AF00",4684=>x"AF00",
4685=>x"AF00",4686=>x"AF00",4687=>x"AF00",4688=>x"AF00",4689=>x"AF00",
4690=>x"AF00",4691=>x"AF00",4692=>x"AF00",4693=>x"AF00",4694=>x"AF00",
4695=>x"AF00",4696=>x"AF00",4697=>x"AF00",4698=>x"AF00",4699=>x"AF00",
4700=>x"AF00",4701=>x"AF00",4702=>x"AF00",4703=>x"AF00",4704=>x"AF00",
4705=>x"AF00",4706=>x"AF00",4707=>x"AF00",4708=>x"AF00",4709=>x"AF00",
4710=>x"AF00",4711=>x"AF00",4712=>x"AF00",4713=>x"AF00",4714=>x"AF00",
4715=>x"AF00",4716=>x"AF00",4717=>x"AF00",4718=>x"AF00",4719=>x"AF00",
4720=>x"AF00",4721=>x"AF00",4722=>x"AF00",4723=>x"AF00",4724=>x"AF00",
4725=>x"AF00",4726=>x"AF00",4727=>x"AF00",4728=>x"AF00",4729=>x"AF00",
4730=>x"AF00",4731=>x"AF00",4732=>x"AF00",4733=>x"AF00",4734=>x"AF00",
4735=>x"AF00",4736=>x"AF00",4737=>x"AF00",4738=>x"AF00",4739=>x"AF00",
4740=>x"AF00",4741=>x"AF00",4742=>x"AF00",4743=>x"AF00",4744=>x"AF00",
4745=>x"AF00",4746=>x"AF00",4747=>x"AF00",4748=>x"AF00",4749=>x"AF00",
4750=>x"AF00",4751=>x"AF00",4752=>x"AF00",4753=>x"AF00",4754=>x"AF00",
4755=>x"AF00",4756=>x"AF00",4757=>x"AF00",4758=>x"AF00",4759=>x"AF00",
4760=>x"AF00",4761=>x"AF00",4762=>x"AF00",4763=>x"AF00",4764=>x"AF00",
4765=>x"AF00",4766=>x"AF00",4767=>x"AF00",4768=>x"AF00",4769=>x"AF00",
4770=>x"AF00",4771=>x"AF00",4772=>x"AF00",4773=>x"AF00",4774=>x"AF00",
4775=>x"AF00",4776=>x"AF00",4777=>x"AF00",4778=>x"AF00",4779=>x"AF00",
4780=>x"AF00",4781=>x"AF00",4782=>x"AF00",4783=>x"AF00",4784=>x"AF00",
4785=>x"AF00",4786=>x"AF00",4787=>x"AF00",4788=>x"AF00",4789=>x"AF00",
4790=>x"AF00",4791=>x"AF00",4792=>x"AF00",4793=>x"AF00",4794=>x"AF00",
4795=>x"AF00",4796=>x"AF00",4797=>x"AF00",4798=>x"AF00",4799=>x"AF00",
4800=>x"AF00",4801=>x"AF00",4802=>x"AF00",4803=>x"AF00",4804=>x"AF00",
4805=>x"AF00",4806=>x"AF00",4807=>x"AF00",4808=>x"AF00",4809=>x"AF00",
4810=>x"AF00",4811=>x"AF00",4812=>x"AF00",4813=>x"AF00",4814=>x"AF00",
4815=>x"AF00",4816=>x"AF00",4817=>x"AF00",4818=>x"AF00",4819=>x"AF00",
4820=>x"AF00",4821=>x"AF00",4822=>x"AF00",4823=>x"AF00",4824=>x"AF00",
4825=>x"AF00",4826=>x"AF00",4827=>x"AF00",4828=>x"AF00",4829=>x"AF00",
4830=>x"AF00",4831=>x"AF00",4832=>x"AF00",4833=>x"AF00",4834=>x"AF00",
4835=>x"AF00",4836=>x"AF00",4837=>x"AF00",4838=>x"AF00",4839=>x"AF00",
4840=>x"AF00",4841=>x"AF00",4842=>x"AF00",4843=>x"AF00",4844=>x"AF00",
4845=>x"AF00",4846=>x"AF00",4847=>x"AF00",4848=>x"AF00",4849=>x"AF00",
4850=>x"AF00",4851=>x"AF00",4852=>x"AF00",4853=>x"AF00",4854=>x"AF00",
4855=>x"AF00",4856=>x"AF00",4857=>x"AF00",4858=>x"AF00",4859=>x"AF00",
4860=>x"AF00",4861=>x"AF00",4862=>x"AF00",4863=>x"AF00",4864=>x"AF00",
4865=>x"AF00",4866=>x"AF00",4867=>x"AF00",4868=>x"AF00",4869=>x"AF00",
4870=>x"AF00",4871=>x"AF00",4872=>x"AF00",4873=>x"AF00",4874=>x"AF00",
4875=>x"AF00",4876=>x"AF00",4877=>x"AF00",4878=>x"AF00",4879=>x"AF00",
4880=>x"AF00",4881=>x"AF00",4882=>x"AF00",4883=>x"AF00",4884=>x"AF00",
4885=>x"AF00",4886=>x"AF00",4887=>x"AF00",4888=>x"AF00",4889=>x"AF00",
4890=>x"AF00",4891=>x"AF00",4892=>x"AF00",4893=>x"AF00",4894=>x"AF00",
4895=>x"AF00",4896=>x"AF00",4897=>x"AF00",4898=>x"AF00",4899=>x"AF00",
4900=>x"AF00",4901=>x"AF00",4902=>x"AF00",4903=>x"AF00",4904=>x"AF00",
4905=>x"AF00",4906=>x"AF00",4907=>x"AF00",4908=>x"AF00",4909=>x"AF00",
4910=>x"AF00",4911=>x"AF00",4912=>x"AF00",4913=>x"AF00",4914=>x"AF00",
4915=>x"AF00",4916=>x"AF00",4917=>x"AF00",4918=>x"AF00",4919=>x"AF00",
4920=>x"AF00",4921=>x"AF00",4922=>x"AF00",4923=>x"AF00",4924=>x"AF00",
4925=>x"AF00",4926=>x"AF00",4927=>x"AF00",4928=>x"AF00",4929=>x"AF00",
4930=>x"AF00",4931=>x"AF00",4932=>x"AF00",4933=>x"AF00",4934=>x"AF00",
4935=>x"AF00",4936=>x"AF00",4937=>x"AF00",4938=>x"AF00",4939=>x"AF00",
4940=>x"AF00",4941=>x"AF00",4942=>x"AF00",4943=>x"AF00",4944=>x"AF00",
4945=>x"AF00",4946=>x"AF00",4947=>x"AF00",4948=>x"AF00",4949=>x"AF00",
4950=>x"AF00",4951=>x"AF00",4952=>x"AF00",4953=>x"AF00",4954=>x"AF00",
4955=>x"AF00",4956=>x"AF00",4957=>x"AF00",4958=>x"AF00",4959=>x"AF00",
4960=>x"AF00",4961=>x"AF00",4962=>x"AF00",4963=>x"AF00",4964=>x"AF00",
4965=>x"AF00",4966=>x"AF00",4967=>x"AF00",4968=>x"AF00",4969=>x"AF00",
4970=>x"AF00",4971=>x"AF00",4972=>x"AF00",4973=>x"AF00",4974=>x"AF00",
4975=>x"AF00",4976=>x"AF00",4977=>x"AF00",4978=>x"AF00",4979=>x"AF00",
4980=>x"AF00",4981=>x"AF00",4982=>x"AF00",4983=>x"AF00",4984=>x"AF00",
4985=>x"AF00",4986=>x"AF00",4987=>x"AF00",4988=>x"AF00",4989=>x"AF00",
4990=>x"AF00",4991=>x"AF00",4992=>x"AF00",4993=>x"AF00",4994=>x"AF00",
4995=>x"AF00",4996=>x"AF00",4997=>x"AF00",4998=>x"AF00",4999=>x"AF00",
5000=>x"AF00",5001=>x"AF00",5002=>x"AF00",5003=>x"AF00",5004=>x"AF00",
5005=>x"AF00",5006=>x"AF00",5007=>x"AF00",5008=>x"AF00",5009=>x"AF00",
5010=>x"AF00",5011=>x"AF00",5012=>x"AF00",5013=>x"AF00",5014=>x"AF00",
5015=>x"AF00",5016=>x"AF00",5017=>x"AF00",5018=>x"AF00",5019=>x"AF00",
5020=>x"AF00",5021=>x"AF00",5022=>x"AF00",5023=>x"AF00",5024=>x"AF00",
5025=>x"AF00",5026=>x"AF00",5027=>x"AF00",5028=>x"AF00",5029=>x"AF00",
5030=>x"AF00",5031=>x"AF00",5032=>x"AF00",5033=>x"AF00",5034=>x"AF00",
5035=>x"AF00",5036=>x"AF00",5037=>x"AF00",5038=>x"AF00",5039=>x"AF00",
5040=>x"AF00",5041=>x"AF00",5042=>x"AF00",5043=>x"AF00",5044=>x"AF00",
5045=>x"AF00",5046=>x"AF00",5047=>x"AF00",5048=>x"AF00",5049=>x"AF00",
5050=>x"AF00",5051=>x"AF00",5052=>x"AF00",5053=>x"AF00",5054=>x"AF00",
5055=>x"AF00",5056=>x"AF00",5057=>x"AF00",5058=>x"AF00",5059=>x"AF00",
5060=>x"AF00",5061=>x"AF00",5062=>x"AF00",5063=>x"AF00",5064=>x"AF00",
5065=>x"AF00",5066=>x"AF00",5067=>x"AF00",5068=>x"AF00",5069=>x"AF00",
5070=>x"AF00",5071=>x"AF00",5072=>x"AF00",5073=>x"AF00",5074=>x"AF00",
5075=>x"AF00",5076=>x"AF00",5077=>x"AF00",5078=>x"AF00",5079=>x"AF00",
5080=>x"AF00",5081=>x"AF00",5082=>x"AF00",5083=>x"AF00",5084=>x"AF00",
5085=>x"AF00",5086=>x"AF00",5087=>x"AF00",5088=>x"AF00",5089=>x"AF00",
5090=>x"AF00",5091=>x"AF00",5092=>x"AF00",5093=>x"AF00",5094=>x"AF00",
5095=>x"AF00",5096=>x"AF00",5097=>x"AF00",5098=>x"AF00",5099=>x"AF00",
5100=>x"AF00",5101=>x"AF00",5102=>x"AF00",5103=>x"AF00",5104=>x"AF00",
5105=>x"AF00",5106=>x"AF00",5107=>x"AF00",5108=>x"AF00",5109=>x"AF00",
5110=>x"AF00",5111=>x"AF00",5112=>x"AF00",5113=>x"AF00",5114=>x"AF00",
5115=>x"AF00",5116=>x"AF00",5117=>x"AF00",5118=>x"AF00",5119=>x"AF00",
5120=>x"AF00",5121=>x"AF00",5122=>x"AF00",5123=>x"AF00",5124=>x"AF00",
5125=>x"AF00",5126=>x"AF00",5127=>x"AF00",5128=>x"AF00",5129=>x"AF00",
5130=>x"AF00",5131=>x"AF00",5132=>x"AF00",5133=>x"AF00",5134=>x"AF00",
5135=>x"AF00",5136=>x"AF00",5137=>x"AF00",5138=>x"AF00",5139=>x"AF00",
5140=>x"AF00",5141=>x"AF00",5142=>x"AF00",5143=>x"AF00",5144=>x"AF00",
5145=>x"AF00",5146=>x"AF00",5147=>x"AF00",5148=>x"AF00",5149=>x"AF00",
5150=>x"AF00",5151=>x"AF00",5152=>x"AF00",5153=>x"AF00",5154=>x"AF00",
5155=>x"AF00",5156=>x"AF00",5157=>x"AF00",5158=>x"AF00",5159=>x"AF00",
5160=>x"AF00",5161=>x"AF00",5162=>x"AF00",5163=>x"AF00",5164=>x"AF00",
5165=>x"AF00",5166=>x"AF00",5167=>x"AF00",5168=>x"AF00",5169=>x"AF00",
5170=>x"AF00",5171=>x"AF00",5172=>x"AF00",5173=>x"AF00",5174=>x"AF00",
5175=>x"AF00",5176=>x"AF00",5177=>x"AF00",5178=>x"AF00",5179=>x"AF00",
5180=>x"AF00",5181=>x"AF00",5182=>x"AF00",5183=>x"AF00",5184=>x"AF00",
5185=>x"AF00",5186=>x"AF00",5187=>x"AF00",5188=>x"AF00",5189=>x"AF00",
5190=>x"AF00",5191=>x"AF00",5192=>x"AF00",5193=>x"AF00",5194=>x"AF00",
5195=>x"AF00",5196=>x"AF00",5197=>x"AF00",5198=>x"AF00",5199=>x"AF00",
5200=>x"AF00",5201=>x"AF00",5202=>x"AF00",5203=>x"AF00",5204=>x"AF00",
5205=>x"AF00",5206=>x"AF00",5207=>x"AF00",5208=>x"AF00",5209=>x"AF00",
5210=>x"AF00",5211=>x"AF00",5212=>x"AF00",5213=>x"AF00",5214=>x"AF00",
5215=>x"AF00",5216=>x"AF00",5217=>x"AF00",5218=>x"AF00",5219=>x"AF00",
5220=>x"AF00",5221=>x"AF00",5222=>x"AF00",5223=>x"AF00",5224=>x"AF00",
5225=>x"AF00",5226=>x"AF00",5227=>x"AF00",5228=>x"AF00",5229=>x"AF00",
5230=>x"AF00",5231=>x"AF00",5232=>x"AF00",5233=>x"AF00",5234=>x"AF00",
5235=>x"AF00",5236=>x"AF00",5237=>x"AF00",5238=>x"AF00",5239=>x"AF00",
5240=>x"AF00",5241=>x"AF00",5242=>x"AF00",5243=>x"AF00",5244=>x"AF00",
5245=>x"AF00",5246=>x"AF00",5247=>x"AF00",5248=>x"AF00",5249=>x"AF00",
5250=>x"AF00",5251=>x"AF00",5252=>x"AF00",5253=>x"AF00",5254=>x"AF00",
5255=>x"AF00",5256=>x"AF00",5257=>x"AF00",5258=>x"AF00",5259=>x"AF00",
5260=>x"AF00",5261=>x"AF00",5262=>x"AF00",5263=>x"AF00",5264=>x"AF00",
5265=>x"AF00",5266=>x"AF00",5267=>x"AF00",5268=>x"AF00",5269=>x"AF00",
5270=>x"AF00",5271=>x"AF00",5272=>x"AF00",5273=>x"AF00",5274=>x"AF00",
5275=>x"AF00",5276=>x"AF00",5277=>x"AF00",5278=>x"AF00",5279=>x"AF00",
5280=>x"AF00",5281=>x"AF00",5282=>x"AF00",5283=>x"AF00",5284=>x"AF00",
5285=>x"AF00",5286=>x"AF00",5287=>x"AF00",5288=>x"AF00",5289=>x"AF00",
5290=>x"AF00",5291=>x"AF00",5292=>x"AF00",5293=>x"AF00",5294=>x"AF00",
5295=>x"AF00",5296=>x"AF00",5297=>x"AF00",5298=>x"AF00",5299=>x"AF00",
5300=>x"AF00",5301=>x"AF00",5302=>x"AF00",5303=>x"AF00",5304=>x"AF00",
5305=>x"AF00",5306=>x"AF00",5307=>x"AF00",5308=>x"AF00",5309=>x"AF00",
5310=>x"AF00",5311=>x"AF00",5312=>x"AF00",5313=>x"AF00",5314=>x"AF00",
5315=>x"AF00",5316=>x"AF00",5317=>x"AF00",5318=>x"AF00",5319=>x"AF00",
5320=>x"AF00",5321=>x"AF00",5322=>x"AF00",5323=>x"AF00",5324=>x"AF00",
5325=>x"AF00",5326=>x"AF00",5327=>x"AF00",5328=>x"AF00",5329=>x"AF00",
5330=>x"AF00",5331=>x"AF00",5332=>x"AF00",5333=>x"AF00",5334=>x"AF00",
5335=>x"AF00",5336=>x"AF00",5337=>x"AF00",5338=>x"AF00",5339=>x"AF00",
5340=>x"AF00",5341=>x"AF00",5342=>x"AF00",5343=>x"AF00",5344=>x"AF00",
5345=>x"AF00",5346=>x"AF00",5347=>x"AF00",5348=>x"AF00",5349=>x"AF00",
5350=>x"AF00",5351=>x"AF00",5352=>x"AF00",5353=>x"AF00",5354=>x"AF00",
5355=>x"AF00",5356=>x"AF00",5357=>x"AF00",5358=>x"AF00",5359=>x"AF00",
5360=>x"AF00",5361=>x"AF00",5362=>x"AF00",5363=>x"AF00",5364=>x"AF00",
5365=>x"AF00",5366=>x"AF00",5367=>x"AF00",5368=>x"AF00",5369=>x"AF00",
5370=>x"AF00",5371=>x"AF00",5372=>x"AF00",5373=>x"AF00",5374=>x"AF00",
5375=>x"AF00",5376=>x"AF00",5377=>x"AF00",5378=>x"AF00",5379=>x"AF00",
5380=>x"AF00",5381=>x"AF00",5382=>x"AF00",5383=>x"AF00",5384=>x"AF00",
5385=>x"AF00",5386=>x"AF00",5387=>x"AF00",5388=>x"AF00",5389=>x"AF00",
5390=>x"AF00",5391=>x"AF00",5392=>x"AF00",5393=>x"AF00",5394=>x"AF00",
5395=>x"AF00",5396=>x"AF00",5397=>x"AF00",5398=>x"AF00",5399=>x"AF00",
5400=>x"AF00",5401=>x"AF00",5402=>x"AF00",5403=>x"AF00",5404=>x"AF00",
5405=>x"AF00",5406=>x"AF00",5407=>x"AF00",5408=>x"AF00",5409=>x"AF00",
5410=>x"AF00",5411=>x"AF00",5412=>x"AF00",5413=>x"AF00",5414=>x"AF00",
5415=>x"AF00",5416=>x"AF00",5417=>x"AF00",5418=>x"AF00",5419=>x"AF00",
5420=>x"AF00",5421=>x"AF00",5422=>x"AF00",5423=>x"AF00",5424=>x"AF00",
5425=>x"AF00",5426=>x"AF00",5427=>x"AF00",5428=>x"AF00",5429=>x"AF00",
5430=>x"AF00",5431=>x"AF00",5432=>x"AF00",5433=>x"AF00",5434=>x"AF00",
5435=>x"AF00",5436=>x"AF00",5437=>x"AF00",5438=>x"AF00",5439=>x"AF00",
5440=>x"AF00",5441=>x"AF00",5442=>x"AF00",5443=>x"AF00",5444=>x"AF00",
5445=>x"AF00",5446=>x"AF00",5447=>x"AF00",5448=>x"AF00",5449=>x"AF00",
5450=>x"AF00",5451=>x"AF00",5452=>x"AF00",5453=>x"AF00",5454=>x"AF00",
5455=>x"AF00",5456=>x"AF00",5457=>x"AF00",5458=>x"AF00",5459=>x"AF00",
5460=>x"AF00",5461=>x"AF00",5462=>x"AF00",5463=>x"AF00",5464=>x"AF00",
5465=>x"AF00",5466=>x"AF00",5467=>x"AF00",5468=>x"AF00",5469=>x"AF00",
5470=>x"AF00",5471=>x"AF00",5472=>x"AF00",5473=>x"AF00",5474=>x"AF00",
5475=>x"AF00",5476=>x"AF00",5477=>x"AF00",5478=>x"AF00",5479=>x"AF00",
5480=>x"AF00",5481=>x"AF00",5482=>x"AF00",5483=>x"AF00",5484=>x"AF00",
5485=>x"AF00",5486=>x"AF00",5487=>x"AF00",5488=>x"AF00",5489=>x"AF00",
5490=>x"AF00",5491=>x"AF00",5492=>x"AF00",5493=>x"AF00",5494=>x"AF00",
5495=>x"AF00",5496=>x"AF00",5497=>x"AF00",5498=>x"AF00",5499=>x"AF00",
5500=>x"AF00",5501=>x"AF00",5502=>x"AF00",5503=>x"AF00",5504=>x"AF00",
5505=>x"AF00",5506=>x"AF00",5507=>x"AF00",5508=>x"AF00",5509=>x"AF00",
5510=>x"AF00",5511=>x"AF00",5512=>x"AF00",5513=>x"AF00",5514=>x"AF00",
5515=>x"AF00",5516=>x"AF00",5517=>x"AF00",5518=>x"AF00",5519=>x"AF00",
5520=>x"AF00",5521=>x"AF00",5522=>x"AF00",5523=>x"AF00",5524=>x"AF00",
5525=>x"AF00",5526=>x"AF00",5527=>x"AF00",5528=>x"AF00",5529=>x"AF00",
5530=>x"AF00",5531=>x"AF00",5532=>x"AF00",5533=>x"AF00",5534=>x"AF00",
5535=>x"AF00",5536=>x"AF00",5537=>x"AF00",5538=>x"AF00",5539=>x"AF00",
5540=>x"AF00",5541=>x"AF00",5542=>x"AF00",5543=>x"AF00",5544=>x"AF00",
5545=>x"AF00",5546=>x"AF00",5547=>x"AF00",5548=>x"AF00",5549=>x"AF00",
5550=>x"AF00",5551=>x"AF00",5552=>x"AF00",5553=>x"AF00",5554=>x"AF00",
5555=>x"AF00",5556=>x"AF00",5557=>x"AF00",5558=>x"AF00",5559=>x"AF00",
5560=>x"AF00",5561=>x"AF00",5562=>x"AF00",5563=>x"AF00",5564=>x"AF00",
5565=>x"AF00",5566=>x"AF00",5567=>x"AF00",5568=>x"AF00",5569=>x"AF00",
5570=>x"AF00",5571=>x"AF00",5572=>x"AF00",5573=>x"AF00",5574=>x"AF00",
5575=>x"AF00",5576=>x"AF00",5577=>x"AF00",5578=>x"AF00",5579=>x"AF00",
5580=>x"AF00",5581=>x"AF00",5582=>x"AF00",5583=>x"AF00",5584=>x"AF00",
5585=>x"AF00",5586=>x"AF00",5587=>x"AF00",5588=>x"AF00",5589=>x"AF00",
5590=>x"AF00",5591=>x"AF00",5592=>x"AF00",5593=>x"AF00",5594=>x"AF00",
5595=>x"AF00",5596=>x"AF00",5597=>x"AF00",5598=>x"AF00",5599=>x"AF00",
5600=>x"AF00",5601=>x"AF00",5602=>x"AF00",5603=>x"AF00",5604=>x"AF00",
5605=>x"AF00",5606=>x"AF00",5607=>x"AF00",5608=>x"AF00",5609=>x"AF00",
5610=>x"AF00",5611=>x"AF00",5612=>x"AF00",5613=>x"AF00",5614=>x"AF00",
5615=>x"AF00",5616=>x"AF00",5617=>x"AF00",5618=>x"AF00",5619=>x"AF00",
5620=>x"AF00",5621=>x"AF00",5622=>x"AF00",5623=>x"AF00",5624=>x"AF00",
5625=>x"AF00",5626=>x"AF00",5627=>x"AF00",5628=>x"AF00",5629=>x"AF00",
5630=>x"AF00",5631=>x"AF00",5632=>x"AF00",5633=>x"AF00",5634=>x"AF00",
5635=>x"AF00",5636=>x"AF00",5637=>x"AF00",5638=>x"AF00",5639=>x"AF00",
5640=>x"AF00",5641=>x"AF00",5642=>x"AF00",5643=>x"AF00",5644=>x"AF00",
5645=>x"AF00",5646=>x"AF00",5647=>x"AF00",5648=>x"AF00",5649=>x"AF00",
5650=>x"AF00",5651=>x"AF00",5652=>x"AF00",5653=>x"AF00",5654=>x"AF00",
5655=>x"AF00",5656=>x"AF00",5657=>x"AF00",5658=>x"AF00",5659=>x"AF00",
5660=>x"AF00",5661=>x"AF00",5662=>x"AF00",5663=>x"AF00",5664=>x"AF00",
5665=>x"AF00",5666=>x"AF00",5667=>x"AF00",5668=>x"AF00",5669=>x"AF00",
5670=>x"AF00",5671=>x"AF00",5672=>x"AF00",5673=>x"AF00",5674=>x"AF00",
5675=>x"AF00",5676=>x"AF00",5677=>x"AF00",5678=>x"AF00",5679=>x"AF00",
5680=>x"AF00",5681=>x"AF00",5682=>x"AF00",5683=>x"AF00",5684=>x"AF00",
5685=>x"AF00",5686=>x"AF00",5687=>x"AF00",5688=>x"AF00",5689=>x"AF00",
5690=>x"AF00",5691=>x"AF00",5692=>x"AF00",5693=>x"AF00",5694=>x"AF00",
5695=>x"AF00",5696=>x"AF00",5697=>x"AF00",5698=>x"AF00",5699=>x"AF00",
5700=>x"AF00",5701=>x"AF00",5702=>x"AF00",5703=>x"AF00",5704=>x"AF00",
5705=>x"AF00",5706=>x"AF00",5707=>x"AF00",5708=>x"AF00",5709=>x"AF00",
5710=>x"AF00",5711=>x"AF00",5712=>x"AF00",5713=>x"AF00",5714=>x"AF00",
5715=>x"AF00",5716=>x"AF00",5717=>x"AF00",5718=>x"AF00",5719=>x"AF00",
5720=>x"AF00",5721=>x"AF00",5722=>x"AF00",5723=>x"AF00",5724=>x"AF00",
5725=>x"AF00",5726=>x"AF00",5727=>x"AF00",5728=>x"AF00",5729=>x"AF00",
5730=>x"AF00",5731=>x"AF00",5732=>x"AF00",5733=>x"AF00",5734=>x"AF00",
5735=>x"AF00",5736=>x"AF00",5737=>x"AF00",5738=>x"AF00",5739=>x"AF00",
5740=>x"AF00",5741=>x"AF00",5742=>x"AF00",5743=>x"AF00",5744=>x"AF00",
5745=>x"AF00",5746=>x"AF00",5747=>x"AF00",5748=>x"AF00",5749=>x"AF00",
5750=>x"AF00",5751=>x"AF00",5752=>x"AF00",5753=>x"AF00",5754=>x"AF00",
5755=>x"AF00",5756=>x"AF00",5757=>x"AF00",5758=>x"AF00",5759=>x"AF00",
5760=>x"AF00",5761=>x"AF00",5762=>x"AF00",5763=>x"AF00",5764=>x"AF00",
5765=>x"AF00",5766=>x"AF00",5767=>x"AF00",5768=>x"AF00",5769=>x"AF00",
5770=>x"AF00",5771=>x"AF00",5772=>x"AF00",5773=>x"AF00",5774=>x"AF00",
5775=>x"AF00",5776=>x"AF00",5777=>x"AF00",5778=>x"AF00",5779=>x"AF00",
5780=>x"AF00",5781=>x"AF00",5782=>x"AF00",5783=>x"AF00",5784=>x"AF00",
5785=>x"AF00",5786=>x"AF00",5787=>x"AF00",5788=>x"AF00",5789=>x"AF00",
5790=>x"AF00",5791=>x"AF00",5792=>x"AF00",5793=>x"AF00",5794=>x"AF00",
5795=>x"AF00",5796=>x"AF00",5797=>x"AF00",5798=>x"AF00",5799=>x"AF00",
5800=>x"AF00",5801=>x"AF00",5802=>x"AF00",5803=>x"AF00",5804=>x"AF00",
5805=>x"AF00",5806=>x"AF00",5807=>x"AF00",5808=>x"AF00",5809=>x"AF00",
5810=>x"AF00",5811=>x"AF00",5812=>x"AF00",5813=>x"AF00",5814=>x"AF00",
5815=>x"AF00",5816=>x"AF00",5817=>x"AF00",5818=>x"AF00",5819=>x"AF00",
5820=>x"AF00",5821=>x"AF00",5822=>x"AF00",5823=>x"AF00",5824=>x"AF00",
5825=>x"AF00",5826=>x"AF00",5827=>x"AF00",5828=>x"AF00",5829=>x"AF00",
5830=>x"AF00",5831=>x"AF00",5832=>x"AF00",5833=>x"AF00",5834=>x"AF00",
5835=>x"AF00",5836=>x"AF00",5837=>x"AF00",5838=>x"AF00",5839=>x"AF00",
5840=>x"AF00",5841=>x"AF00",5842=>x"AF00",5843=>x"AF00",5844=>x"AF00",
5845=>x"AF00",5846=>x"AF00",5847=>x"AF00",5848=>x"AF00",5849=>x"AF00",
5850=>x"AF00",5851=>x"AF00",5852=>x"AF00",5853=>x"AF00",5854=>x"AF00",
5855=>x"AF00",5856=>x"AF00",5857=>x"AF00",5858=>x"AF00",5859=>x"AF00",
5860=>x"AF00",5861=>x"AF00",5862=>x"AF00",5863=>x"AF00",5864=>x"AF00",
5865=>x"AF00",5866=>x"AF00",5867=>x"AF00",5868=>x"AF00",5869=>x"AF00",
5870=>x"AF00",5871=>x"AF00",5872=>x"AF00",5873=>x"AF00",5874=>x"AF00",
5875=>x"AF00",5876=>x"AF00",5877=>x"AF00",5878=>x"AF00",5879=>x"AF00",
5880=>x"AF00",5881=>x"AF00",5882=>x"AF00",5883=>x"AF00",5884=>x"AF00",
5885=>x"AF00",5886=>x"AF00",5887=>x"AF00",5888=>x"AF00",5889=>x"AF00",
5890=>x"AF00",5891=>x"AF00",5892=>x"AF00",5893=>x"AF00",5894=>x"AF00",
5895=>x"AF00",5896=>x"AF00",5897=>x"AF00",5898=>x"AF00",5899=>x"AF00",
5900=>x"AF00",5901=>x"AF00",5902=>x"AF00",5903=>x"AF00",5904=>x"AF00",
5905=>x"AF00",5906=>x"AF00",5907=>x"AF00",5908=>x"AF00",5909=>x"AF00",
5910=>x"AF00",5911=>x"AF00",5912=>x"AF00",5913=>x"AF00",5914=>x"AF00",
5915=>x"AF00",5916=>x"AF00",5917=>x"AF00",5918=>x"AF00",5919=>x"AF00",
5920=>x"AF00",5921=>x"AF00",5922=>x"AF00",5923=>x"AF00",5924=>x"AF00",
5925=>x"AF00",5926=>x"AF00",5927=>x"AF00",5928=>x"AF00",5929=>x"AF00",
5930=>x"AF00",5931=>x"AF00",5932=>x"AF00",5933=>x"AF00",5934=>x"AF00",
5935=>x"AF00",5936=>x"AF00",5937=>x"AF00",5938=>x"AF00",5939=>x"AF00",
5940=>x"AF00",5941=>x"AF00",5942=>x"AF00",5943=>x"AF00",5944=>x"AF00",
5945=>x"AF00",5946=>x"AF00",5947=>x"AF00",5948=>x"AF00",5949=>x"AF00",
5950=>x"AF00",5951=>x"AF00",5952=>x"AF00",5953=>x"AF00",5954=>x"AF00",
5955=>x"AF00",5956=>x"AF00",5957=>x"AF00",5958=>x"AF00",5959=>x"AF00",
5960=>x"AF00",5961=>x"AF00",5962=>x"AF00",5963=>x"AF00",5964=>x"AF00",
5965=>x"AF00",5966=>x"AF00",5967=>x"AF00",5968=>x"AF00",5969=>x"AF00",
5970=>x"AF00",5971=>x"AF00",5972=>x"AF00",5973=>x"AF00",5974=>x"AF00",
5975=>x"AF00",5976=>x"AF00",5977=>x"AF00",5978=>x"AF00",5979=>x"AF00",
5980=>x"AF00",5981=>x"AF00",5982=>x"AF00",5983=>x"AF00",5984=>x"AF00",
5985=>x"AF00",5986=>x"AF00",5987=>x"AF00",5988=>x"AF00",5989=>x"AF00",
5990=>x"AF00",5991=>x"AF00",5992=>x"AF00",5993=>x"AF00",5994=>x"AF00",
5995=>x"AF00",5996=>x"AF00",5997=>x"AF00",5998=>x"AF00",5999=>x"AF00",
6000=>x"AF00",6001=>x"AF00",6002=>x"AF00",6003=>x"AF00",6004=>x"AF00",
6005=>x"AF00",6006=>x"AF00",6007=>x"AF00",6008=>x"AF00",6009=>x"AF00",
6010=>x"AF00",6011=>x"AF00",6012=>x"AF00",6013=>x"AF00",6014=>x"AF00",
6015=>x"AF00",6016=>x"AF00",6017=>x"AF00",6018=>x"AF00",6019=>x"AF00",
6020=>x"AF00",6021=>x"AF00",6022=>x"AF00",6023=>x"AF00",6024=>x"AF00",
6025=>x"AF00",6026=>x"AF00",6027=>x"AF00",6028=>x"AF00",6029=>x"AF00",
6030=>x"AF00",6031=>x"AF00",6032=>x"AF00",6033=>x"AF00",6034=>x"AF00",
6035=>x"AF00",6036=>x"AF00",6037=>x"AF00",6038=>x"AF00",6039=>x"AF00",
6040=>x"AF00",6041=>x"AF00",6042=>x"AF00",6043=>x"AF00",6044=>x"AF00",
6045=>x"AF00",6046=>x"AF00",6047=>x"AF00",6048=>x"AF00",6049=>x"AF00",
6050=>x"AF00",6051=>x"AF00",6052=>x"AF00",6053=>x"AF00",6054=>x"AF00",
6055=>x"AF00",6056=>x"AF00",6057=>x"AF00",6058=>x"AF00",6059=>x"AF00",
6060=>x"AF00",6061=>x"AF00",6062=>x"AF00",6063=>x"AF00",6064=>x"AF00",
6065=>x"AF00",6066=>x"AF00",6067=>x"AF00",6068=>x"AF00",6069=>x"AF00",
6070=>x"AF00",6071=>x"AF00",6072=>x"AF00",6073=>x"AF00",6074=>x"AF00",
6075=>x"AF00",6076=>x"AF00",6077=>x"AF00",6078=>x"AF00",6079=>x"AF00",
6080=>x"AF00",6081=>x"AF00",6082=>x"AF00",6083=>x"AF00",6084=>x"AF00",
6085=>x"AF00",6086=>x"AF00",6087=>x"AF00",6088=>x"AF00",6089=>x"AF00",
6090=>x"AF00",6091=>x"AF00",6092=>x"AF00",6093=>x"AF00",6094=>x"AF00",
6095=>x"AF00",6096=>x"AF00",6097=>x"AF00",6098=>x"AF00",6099=>x"AF00",
6100=>x"AF00",6101=>x"AF00",6102=>x"AF00",6103=>x"AF00",6104=>x"AF00",
6105=>x"AF00",6106=>x"AF00",6107=>x"AF00",6108=>x"AF00",6109=>x"AF00",
6110=>x"AF00",6111=>x"AF00",6112=>x"AF00",6113=>x"AF00",6114=>x"AF00",
6115=>x"AF00",6116=>x"AF00",6117=>x"AF00",6118=>x"AF00",6119=>x"AF00",
6120=>x"AF00",6121=>x"AF00",6122=>x"AF00",6123=>x"AF00",6124=>x"AF00",
6125=>x"AF00",6126=>x"AF00",6127=>x"AF00",6128=>x"AF00",6129=>x"AF00",
6130=>x"AF00",6131=>x"AF00",6132=>x"AF00",6133=>x"AF00",6134=>x"AF00",
6135=>x"AF00",6136=>x"AF00",6137=>x"AF00",6138=>x"AF00",6139=>x"AF00",
OTHERS => x"0000"
);
BEGIN
	data <= ram(to_uint(addr)) WHEN re
	   ELSE x"ZZZZ";
	
	PROCESS(ALL) IS BEGIN
		IF rising_edge(clk) THEN
		IF NOT re AND we THEN
			ram(to_uint(addr)) <= data;
		END IF;
		END IF;
	END PROCESS;
	

END ARCHITECTURE arch;

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY Gowin_rPLL IS
	PORT(
		clkout :   OUT std_ulogic;
		clkin  : IN    std_ulogic
	);
END ENTITY Gowin_rPLL;

ARCHITECTURE Behavioral OF Gowin_rPLL IS
BEGIN
	clkout <= clkin;
END ARCHITECTURE;
